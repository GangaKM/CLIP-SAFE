magic
tech sky130A
magscale 1 2
timestamp 1698651669
<< pwell >>
rect 644 1146 681 1291
rect 1630 1192 1660 1286
<< locali >>
rect 223 2021 3623 2056
rect 223 1919 3623 1979
rect 1279 1810 1347 1919
rect 2435 1812 2503 1919
rect 1101 1688 1524 1725
rect 2262 1689 2685 1726
rect 1132 1172 1549 1215
rect 2287 1199 2706 1208
rect 2287 1166 2707 1199
rect 1301 998 1376 1096
rect 2464 998 2532 1100
rect 226 932 3625 998
rect 3624 890 3625 932
rect 226 860 3625 890
rect 2748 478 2932 628
<< viali >>
rect 218 1979 3627 2021
rect 215 890 3624 932
<< metal1 >>
rect 206 2021 3639 2027
rect 206 1979 218 2021
rect 3627 1979 3639 2021
rect 206 1973 3639 1979
rect 206 1916 3616 1973
rect 206 1195 248 1916
rect 418 1675 428 1742
rect 483 1675 493 1742
rect 604 1716 681 1753
rect 604 1708 641 1716
rect 642 1708 681 1716
rect 604 1671 681 1708
rect 642 1636 681 1671
rect 804 1668 814 1735
rect 869 1668 879 1735
rect 988 1666 1066 1753
rect 1589 1676 1621 1916
rect 1670 1807 2115 1850
rect 541 1279 570 1632
rect 644 1441 681 1636
rect 904 1580 914 1632
rect 976 1580 986 1632
rect 1033 1442 1066 1666
rect 1759 1665 1842 1702
rect 1805 1629 1842 1665
rect 1719 1576 1844 1629
rect 1033 1441 1744 1442
rect 642 1411 1744 1441
rect 444 1195 454 1203
rect 206 1153 454 1195
rect 444 1136 454 1153
rect 509 1136 519 1203
rect 644 1146 681 1411
rect 1033 1409 1744 1411
rect 915 1269 925 1321
rect 987 1269 997 1321
rect 836 1133 846 1200
rect 901 1133 911 1200
rect 1033 1145 1066 1409
rect 1600 1134 1610 1194
rect 1666 1134 1676 1194
rect 302 1061 597 1100
rect 1711 1064 1744 1409
rect 1805 1146 1842 1576
rect 1973 1241 2007 1762
rect 2161 1679 2193 1916
rect 2743 1759 2776 1770
rect 2743 1659 2784 1759
rect 2907 1665 2917 1732
rect 2972 1665 2982 1732
rect 2743 1442 2776 1659
rect 2814 1576 2824 1628
rect 2889 1576 2899 1628
rect 2099 1440 2776 1442
rect 3118 1440 3155 1761
rect 3295 1673 3305 1740
rect 3360 1673 3370 1740
rect 2099 1410 3155 1440
rect 2099 1409 2776 1410
rect 1973 1162 2046 1241
rect 2099 1068 2132 1409
rect 2743 1240 2776 1409
rect 2842 1268 2852 1320
rect 2917 1268 2927 1320
rect 2164 1139 2174 1199
rect 2229 1139 2239 1199
rect 2743 1143 2818 1240
rect 3118 1239 3155 1410
rect 3238 1273 3278 1621
rect 2939 1147 2949 1214
rect 3004 1147 3014 1214
rect 3118 1128 3198 1239
rect 3324 1147 3334 1214
rect 3389 1195 3399 1214
rect 3389 1193 3429 1195
rect 3562 1193 3602 1916
rect 3389 1154 3602 1193
rect 3389 1153 3528 1154
rect 3389 1147 3399 1153
rect 3240 1096 3528 1101
rect 2878 1064 3528 1096
rect 2878 1058 3311 1064
rect 280 956 290 997
rect 223 940 290 956
rect 361 956 371 997
rect 3474 956 3484 1001
rect 361 940 3484 956
rect 223 938 3484 940
rect 203 932 3484 938
rect 3541 956 3551 1001
rect 3541 938 3626 956
rect 3541 932 3636 938
rect 203 890 215 932
rect 3624 890 3636 932
rect 203 884 3636 890
rect 223 853 3626 884
rect 2740 750 2750 808
rect 2932 750 2942 808
<< via1 >>
rect 428 1675 483 1742
rect 814 1668 869 1735
rect 914 1580 976 1632
rect 454 1136 509 1203
rect 925 1269 987 1321
rect 846 1133 901 1200
rect 1610 1134 1666 1194
rect 2917 1665 2972 1732
rect 2824 1576 2889 1628
rect 3305 1673 3360 1740
rect 2852 1268 2917 1320
rect 2174 1139 2229 1199
rect 2949 1147 3004 1214
rect 3334 1147 3389 1214
rect 290 940 361 997
rect 3484 932 3541 1001
rect 2750 750 2932 808
<< metal2 >>
rect 919 1845 949 1860
rect 880 1814 965 1845
rect 428 1742 483 1752
rect 385 1739 428 1740
rect 306 1696 428 1739
rect 306 1007 349 1696
rect 385 1695 428 1696
rect 409 1691 428 1695
rect 814 1735 869 1745
rect 483 1691 814 1727
rect 428 1665 483 1675
rect 814 1658 869 1668
rect 919 1642 949 1814
rect 2917 1732 2972 1742
rect 3305 1740 3360 1750
rect 2972 1682 3305 1718
rect 2917 1655 2972 1665
rect 3360 1676 3526 1718
rect 3305 1663 3360 1673
rect 914 1632 976 1642
rect 914 1570 976 1580
rect 2824 1630 2889 1638
rect 2824 1628 2890 1630
rect 2889 1576 2890 1628
rect 922 1331 957 1570
rect 2824 1566 2890 1576
rect 1630 1371 2209 1401
rect 922 1321 987 1331
rect 922 1278 925 1321
rect 925 1259 987 1269
rect 454 1203 509 1213
rect 439 1143 454 1179
rect 846 1200 901 1210
rect 1630 1204 1660 1371
rect 2179 1209 2209 1371
rect 2854 1330 2890 1566
rect 2852 1320 2917 1330
rect 2852 1258 2917 1268
rect 2949 1214 3004 1224
rect 509 1143 846 1179
rect 454 1126 509 1136
rect 846 1123 901 1133
rect 1610 1194 1666 1204
rect 1610 1124 1666 1134
rect 2174 1199 2229 1209
rect 2229 1152 2810 1192
rect 2944 1157 2949 1193
rect 2174 1129 2229 1139
rect 290 997 361 1007
rect 290 930 361 940
rect 2770 826 2810 1152
rect 3334 1214 3389 1224
rect 3004 1157 3334 1193
rect 2949 1137 3004 1147
rect 3389 1157 3395 1193
rect 3334 1137 3389 1147
rect 3484 1011 3526 1676
rect 3484 1001 3541 1011
rect 3484 922 3541 932
rect 2750 808 2946 826
rect 2736 764 2750 793
rect 2932 750 2946 808
rect 2750 740 2932 750
use sky130_fd_pr__nfet_01v8_SMGLWN  XM1
timestamp 1698155087
transform 1 0 1340 0 1 1186
box -246 -260 246 260
use sky130_fd_pr__nfet_01v8_SMGLWN  XM2
timestamp 1698155087
transform 1 0 2498 0 1 1186
box -246 -260 246 260
use sky130_fd_pr__pfet_01v8_TM5SY6  XM3
timestamp 1698155087
transform 1 0 1313 0 1 1716
box -246 -269 246 269
use sky130_fd_pr__pfet_01v8_TM5SY6  XM4
timestamp 1698155087
transform 1 0 541 0 1 1716
box -246 -269 246 269
use sky130_fd_pr__pfet_01v8_TM5SY6  XM5
timestamp 1698155087
transform 1 0 1699 0 1 1716
box -246 -269 246 269
use sky130_fd_pr__pfet_01v8_TM5SY6  XM6
timestamp 1698155087
transform 1 0 2085 0 1 1716
box -246 -269 246 269
use sky130_fd_pr__nfet_01v8_SMGLWN  XM7
timestamp 1698155087
transform 1 0 1726 0 1 1186
box -246 -260 246 260
use sky130_fd_pr__nfet_01v8_SMGLWN  XM8
timestamp 1698155087
transform 1 0 2112 0 1 1186
box -246 -260 246 260
use sky130_fd_pr__nfet_01v8_PVEW3M  XM9
timestamp 1697998059
transform 0 1 2839 -1 0 685
box -246 -310 246 310
use sky130_fd_pr__nfet_01v8_SMGLWN  XM10
timestamp 1698155087
transform 1 0 568 0 1 1186
box -246 -260 246 260
use sky130_fd_pr__nfet_01v8_SMGLWN  XM11
timestamp 1698155087
transform 1 0 954 0 1 1186
box -246 -260 246 260
use sky130_fd_pr__pfet_01v8_TM5SY6  XM12
timestamp 1698155087
transform 1 0 927 0 1 1716
box -246 -269 246 269
use sky130_fd_pr__nfet_01v8_SMGLWN  XM13
timestamp 1698155087
transform 1 0 2884 0 1 1186
box -246 -260 246 260
use sky130_fd_pr__nfet_01v8_SMGLWN  XM14
timestamp 1698155087
transform 1 0 3270 0 1 1186
box -246 -260 246 260
use sky130_fd_pr__pfet_01v8_TM5SY6  XM15
timestamp 1698155087
transform 1 0 2857 0 1 1716
box -246 -269 246 269
use sky130_fd_pr__pfet_01v8_TM5SY6  XM16
timestamp 1698155087
transform 1 0 3243 0 1 1716
box -246 -269 246 269
use sky130_fd_pr__pfet_01v8_TM5SY6  XM18
timestamp 1698155087
transform 1 0 2471 0 1 1716
box -246 -269 246 269
<< labels >>
rlabel locali 1990 2056 1990 2056 1 Vdd
rlabel metal1 2801 1440 2801 1440 1 Vcm
rlabel metal1 1405 853 1405 853 5 gnd
<< end >>
