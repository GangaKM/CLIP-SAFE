magic
tech sky130A
magscale 1 2
timestamp 1698849032
<< nwell >>
rect 6148 -686 12052 -44
rect 13860 -744 14344 -470
rect 17266 -622 25072 -74
<< nsubdiff >>
rect 13966 -536 14244 -508
rect 13966 -680 14002 -536
rect 14210 -680 14244 -536
rect 13966 -704 14244 -680
<< nsubdiffcont >>
rect 14002 -680 14210 -536
<< locali >>
rect 13966 -536 14244 -508
rect 13966 -680 14002 -536
rect 14210 -680 14244 -536
rect 13966 -704 14244 -680
<< viali >>
rect 14002 -680 14210 -536
<< metal1 >>
rect 6228 9446 7456 9628
rect 3840 7248 4258 8522
rect 3840 7072 4226 7248
rect 3718 7056 4226 7072
rect 3710 6990 4226 7056
rect 3710 6338 3780 6990
rect 4114 6338 4226 6990
rect 3710 6278 4226 6338
rect 3718 6274 4226 6278
rect 3840 1124 4226 6274
rect 4490 6886 4930 6982
rect 4490 6012 4592 6886
rect 4850 6012 4930 6886
rect 4490 5952 4930 6012
rect 3840 -274 4306 1124
rect 4558 94 4916 5952
rect 26076 3850 26578 5842
rect 25236 3740 25668 3806
rect 25236 3272 25360 3740
rect 25600 3272 25668 3740
rect 4558 -146 12752 94
rect 25236 92 25668 3272
rect 26076 3344 26160 3850
rect 26492 3590 26578 3850
rect 26492 3344 26576 3590
rect 26076 3266 26576 3344
rect 26100 2984 26506 3266
rect 25918 186 26506 2984
rect 13472 -10 14786 58
rect 13472 -42 13532 -10
rect 3840 -1238 4226 -274
rect 4582 -338 12752 -146
rect 13460 -300 13532 -42
rect 14726 -300 14786 -10
rect 13460 -380 14786 -300
rect 16204 -340 25668 92
rect 13460 -480 14774 -380
rect 13996 -508 14202 -480
rect 13966 -536 14244 -508
rect 5062 -1226 6078 -548
rect 13966 -680 14002 -536
rect 14210 -680 14244 -536
rect 13966 -704 14244 -680
rect 14922 -622 15628 -556
rect 14922 -832 15012 -622
rect 13863 -865 14216 -832
rect 14868 -836 15012 -832
rect 14748 -869 15012 -836
rect 14868 -873 15012 -869
rect 14922 -878 15012 -873
rect 15478 -878 15628 -622
rect 14922 -950 15628 -878
rect 13488 -1052 13522 -978
rect 13706 -1052 13740 -978
rect 14384 -1040 14418 -982
rect 14602 -1040 14636 -982
rect 13954 -1052 14212 -1046
rect 14380 -1052 14418 -1040
rect 14598 -1052 14636 -1040
rect 13452 -1120 14688 -1052
rect 4354 -1238 12656 -1226
rect 3840 -1542 12656 -1238
rect 3910 -1634 12656 -1542
rect 13452 -1494 13558 -1120
rect 14540 -1494 14688 -1120
rect 16470 -1154 25128 -544
rect 26100 -1154 26506 186
rect 16470 -1178 26506 -1154
rect 13452 -1566 14688 -1494
rect 16012 -1562 26506 -1178
rect 16012 -1610 26386 -1562
rect 5062 -1646 6078 -1634
rect 25068 -1658 26386 -1610
<< via1 >>
rect 3780 6338 4114 6990
rect 4592 6012 4850 6886
rect 25360 3272 25600 3740
rect 26160 3344 26492 3850
rect 13532 -300 14726 -10
rect 15012 -878 15478 -622
rect 13558 -1494 14540 -1120
<< metal2 >>
rect 3718 6990 4214 7072
rect 3718 6338 3780 6990
rect 4114 6338 4214 6990
rect 3718 6274 4214 6338
rect 4490 6886 4930 6982
rect 4490 6012 4592 6886
rect 4850 6012 4930 6886
rect 4490 5952 4930 6012
rect 26076 3850 26576 3934
rect 25250 3740 25666 3792
rect 25250 3272 25360 3740
rect 25600 3272 25666 3740
rect 25250 3206 25666 3272
rect 26076 3344 26160 3850
rect 26492 3344 26576 3850
rect 26076 3266 26576 3344
rect 13472 -10 14786 58
rect 13472 -300 13532 -10
rect 14726 -300 14786 -10
rect 13472 -380 14786 -300
rect 12638 -612 13352 -546
rect 12638 -878 12738 -612
rect 13226 -878 13352 -612
rect 12638 -930 13352 -878
rect 14922 -622 15628 -556
rect 14922 -878 15012 -622
rect 15478 -878 15628 -622
rect 14922 -950 15628 -878
rect 13452 -1120 14688 -1052
rect 13452 -1494 13558 -1120
rect 14540 -1494 14688 -1120
rect 13452 -1566 14688 -1494
<< via2 >>
rect 3780 6338 4114 6990
rect 4592 6012 4850 6886
rect 25360 3272 25600 3740
rect 26160 3344 26492 3850
rect 13532 -300 14726 -10
rect 12738 -878 13226 -612
rect 15012 -878 15478 -622
rect 13558 -1494 14540 -1120
<< metal3 >>
rect 3718 6990 4214 7072
rect 3718 6338 3780 6990
rect 4114 6338 4214 6990
rect 3718 6274 4214 6338
rect 4490 6886 4930 6982
rect 4490 6012 4592 6886
rect 4850 6012 4930 6886
rect 4490 5952 4930 6012
rect 26076 3850 26576 3934
rect 25250 3740 25666 3792
rect 25250 3272 25360 3740
rect 25600 3272 25666 3740
rect 25250 3206 25666 3272
rect 26076 3344 26160 3850
rect 26492 3344 26576 3850
rect 26076 3266 26576 3344
rect 13472 -10 14786 58
rect 13472 -300 13532 -10
rect 14726 -300 14786 -10
rect 13472 -380 14786 -300
rect 4960 -546 13254 -538
rect 4960 -612 13352 -546
rect 15476 -556 15562 1695
rect 4960 -878 12738 -612
rect 13226 -878 13352 -612
rect 4960 -930 13352 -878
rect 14922 -622 26624 -556
rect 14922 -878 15012 -622
rect 15478 -878 26624 -622
rect 14922 -948 26624 -878
rect 14922 -950 15628 -948
rect 13452 -1120 14688 -1052
rect 13452 -1494 13558 -1120
rect 14540 -1494 14688 -1120
rect 13452 -1566 14688 -1494
<< via3 >>
rect 3780 6338 4114 6990
rect 4592 6012 4850 6886
rect 25360 3272 25600 3740
rect 26160 3344 26492 3850
rect 13532 -300 14726 -10
rect 13558 -1494 14540 -1120
<< metal4 >>
rect 3718 6990 4214 7072
rect 3718 6338 3780 6990
rect 4114 6338 4214 6990
rect 3718 6274 4214 6338
rect 4314 227 4972 5569
rect 25147 3740 25845 8873
rect 25147 3272 25360 3740
rect 25600 3272 25845 3740
rect 25147 227 25845 3272
rect 26076 3850 26576 3934
rect 26076 3344 26160 3850
rect 26492 3344 26576 3850
rect 26076 3266 26576 3344
rect 4313 -10 26624 227
rect 4313 -300 13532 -10
rect 14726 -300 26624 -10
rect 4313 -471 26624 -300
rect 13452 -1120 14688 -1052
rect 13452 -1494 13558 -1120
rect 14540 -1494 14688 -1120
rect 13452 -1566 14688 -1494
<< via4 >>
rect 3780 6344 4108 6986
rect 26160 3344 26492 3850
rect 13558 -1494 14540 -1120
<< metal5 >>
rect 3739 10192 4397 10505
rect 3720 6986 4397 10192
rect 3720 6344 3780 6986
rect 4108 6344 4397 6986
rect 3720 -1049 4397 6344
rect 25999 3850 26589 4745
rect 25999 3344 26160 3850
rect 26492 3344 26589 3850
rect 3720 -1088 25272 -1049
rect 25999 -1088 26589 3344
rect 3720 -1120 26624 -1088
rect 3720 -1494 13558 -1120
rect 14540 -1494 26624 -1120
rect 3720 -1707 26624 -1494
rect 3739 -1767 26624 -1707
rect 25999 -1785 26589 -1767
use buffer_digital  buffer_digital_0 ~/Desktop/charge_pumps2/layout_files
timestamp 1698771642
transform 1 0 14386 0 1 -1016
box -274 0 415 576
use buffer_digital  buffer_digital_1
timestamp 1698771642
transform 1 0 13490 0 1 -1012
box -274 0 415 576
use charge_pump  charge_pump_0 ~/Desktop/charge_pumps2/layout_files2
timestamp 1698849032
transform 1 0 2956 0 1 9440
box 764 -7862 23794 19014
use nmos_decap_10  nmos_decap_10_0
timestamp 1698837560
transform 0 1 4166 -1 0 842
box -10 -42 1060 416
use nmos_decap_10  nmos_decap_10_1
timestamp 1698837560
transform 0 1 4166 -1 0 1802
box -10 -42 1060 416
use nmos_decap_10  nmos_decap_10_2
timestamp 1698837560
transform 0 1 4166 -1 0 2762
box -10 -42 1060 416
use nmos_decap_10  nmos_decap_10_3
timestamp 1698837560
transform 0 1 4166 -1 0 3722
box -10 -42 1060 416
use nmos_decap_10  nmos_decap_10_4
timestamp 1698837560
transform 0 1 4166 -1 0 4682
box -10 -42 1060 416
use nmos_decap_10  nmos_decap_10_5
timestamp 1698837560
transform 0 1 4166 -1 0 5642
box -10 -42 1060 416
use nmos_decap_10  nmos_decap_10_6
timestamp 1698837560
transform 0 1 25530 1 0 190
box -10 -42 1060 416
use nmos_decap_10  nmos_decap_10_7
timestamp 1698837560
transform 0 1 25530 1 0 1150
box -10 -42 1060 416
use nmos_decap_10  nmos_decap_10_8
timestamp 1698837560
transform 0 1 25530 1 0 2110
box -10 -42 1060 416
use pmos_decap_10  pmos_decap_10_0
timestamp 1698841269
transform 1 0 5194 0 -1 -206
box 0 -108 1098 464
use pmos_decap_10  pmos_decap_10_1
timestamp 1698841269
transform 1 0 6266 0 -1 -196
box 0 -108 1098 464
use pmos_decap_10  pmos_decap_10_2
timestamp 1698841269
transform 1 0 7338 0 -1 -174
box 0 -108 1098 464
use pmos_decap_10  pmos_decap_10_3
timestamp 1698841269
transform 1 0 8410 0 -1 -178
box 0 -108 1098 464
use pmos_decap_10  pmos_decap_10_4
timestamp 1698841269
transform 1 0 9482 0 -1 -178
box 0 -108 1098 464
use pmos_decap_10  pmos_decap_10_5
timestamp 1698841269
transform 1 0 10554 0 -1 -178
box 0 -108 1098 464
use pmos_decap_10  pmos_decap_10_6
timestamp 1698841269
transform 1 0 16414 0 -1 -186
box 0 -108 1098 464
use pmos_decap_10  pmos_decap_10_7
timestamp 1698841269
transform 1 0 17486 0 -1 -182
box 0 -108 1098 464
use pmos_decap_10  pmos_decap_10_8
timestamp 1698841269
transform 1 0 18558 0 -1 -176
box 0 -108 1098 464
use pmos_decap_10  pmos_decap_10_9
timestamp 1698841269
transform 1 0 19630 0 -1 -174
box 0 -108 1098 464
use pmos_decap_10  pmos_decap_10_10
timestamp 1698841269
transform 1 0 20702 0 -1 -174
box 0 -108 1098 464
use pmos_decap_10  pmos_decap_10_11
timestamp 1698841269
transform 1 0 21774 0 -1 -174
box 0 -108 1098 464
use pmos_decap_10  pmos_decap_10_12
timestamp 1698841269
transform 1 0 22846 0 -1 -180
box 0 -108 1098 464
use pmos_decap_10  pmos_decap_10_13
timestamp 1698841269
transform 1 0 23918 0 -1 -176
box 0 -108 1098 464
<< end >>
