* SPICE3 file created from comparator_final_compact.ext - technology: sky130A

.subckt sky130_fd_pr__nfet_01v8_GWFSUW a_15_n130# a_63_n42# a_n177_n130# a_255_n42#
+ a_n129_n42# a_111_64# a_n321_n42# a_159_n42# a_n81_64# a_n273_64# a_351_n42# a_207_n130#
+ a_303_64# a_n33_n42# a_n369_n130# a_n225_n42# a_n413_n42# VSUBS
X0 a_63_n42# a_15_n130# a_n33_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X1 a_n33_n42# a_n81_64# a_n129_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X2 a_351_n42# a_303_64# a_255_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X3 a_159_n42# a_111_64# a_63_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X4 a_255_n42# a_207_n130# a_159_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X5 a_n321_n42# a_n369_n130# a_n413_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X6 a_n225_n42# a_n273_64# a_n321_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X7 a_n129_n42# a_n177_n130# a_n225_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
.ends

.subckt sky130_fd_pr__pfet_01v8_BH9SS5 w_n246_n319# a_n50_n197# a_50_n100# a_n108_n100#
+ VSUBS
X0 a_50_n100# a_n50_n197# a_n108_n100# w_n246_n319# sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
.ends

.subckt sky130_fd_pr__nfet_01v8_53744R a_n210_n274# a_50_n100# a_n108_n100# a_n50_n188#
X0 a_50_n100# a_n50_n188# a_n108_n100# a_n210_n274# sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
.ends

.subckt inverter m1_176_134# m1_272_214# li_n18_880# VSUBS
Xsky130_fd_pr__pfet_01v8_BH9SS5_0 li_n18_880# m1_176_134# m1_272_214# li_n18_880#
+ VSUBS sky130_fd_pr__pfet_01v8_BH9SS5
Xsky130_fd_pr__nfet_01v8_53744R_0 VSUBS m1_272_214# VSUBS m1_176_134# sky130_fd_pr__nfet_01v8_53744R
.ends

.subckt sky130_fd_pr__nfet_01v8_PVEW3M a_n210_n274# a_50_n100# a_n108_n100# a_n50_n188#
X0 a_50_n100# a_n50_n188# a_n108_n100# a_n210_n274# sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
.ends

.subckt sky130_fd_pr__pfet_01v8_X3YSY6 w_n246_n319# a_n50_n197# a_50_n100# a_n108_n100#
+ VSUBS
X0 a_50_n100# a_n50_n197# a_n108_n100# w_n246_n319# sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
.ends

.subckt sky130_fd_pr__pfet_01v8_B5E2Q5 w_n246_n319# a_n50_n197# a_50_n100# a_n108_n100#
+ VSUBS
X0 a_50_n100# a_n50_n197# a_n108_n100# w_n246_n319# sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
.ends

.subckt comparator_layout m1_1704_1482# m1_1411_1896# m1_2488_2128# li_905_2237# m1_2014_1251#
+ XM33/a_n50_n188# XM34/a_n50_n188# m1_1061_1257# m1_852_1342# VSUBS XM25/a_n50_n188#
+ XM26/a_n50_n188#
XXM34 VSUBS m1_852_1342# m1_2014_1251# XM34/a_n50_n188# sky130_fd_pr__nfet_01v8_PVEW3M
XXM35 VSUBS VSUBS m1_852_1342# m1_2488_2128# sky130_fd_pr__nfet_01v8_PVEW3M
XXM25 VSUBS m1_1061_1257# m1_852_1342# XM25/a_n50_n188# sky130_fd_pr__nfet_01v8_PVEW3M
XXM26 VSUBS m1_1061_1257# m1_852_1342# XM26/a_n50_n188# sky130_fd_pr__nfet_01v8_PVEW3M
XXM27 VSUBS m1_1411_1896# m1_1061_1257# m1_1704_1482# sky130_fd_pr__nfet_01v8_PVEW3M
XXM28 VSUBS m1_1704_1482# m1_2014_1251# m1_1411_1896# sky130_fd_pr__nfet_01v8_PVEW3M
XXM29 li_905_2237# m1_2488_2128# m1_1411_1896# li_905_2237# VSUBS sky130_fd_pr__pfet_01v8_X3YSY6
Xsky130_fd_pr__pfet_01v8_B5E2Q5_0 li_905_2237# m1_2488_2128# m1_2014_1251# m1_1061_1257#
+ VSUBS sky130_fd_pr__pfet_01v8_B5E2Q5
XXM30 li_905_2237# m1_1704_1482# m1_1411_1896# li_905_2237# VSUBS sky130_fd_pr__pfet_01v8_X3YSY6
XXM31 li_905_2237# m1_1411_1896# m1_1704_1482# li_905_2237# VSUBS sky130_fd_pr__pfet_01v8_X3YSY6
XXM32 li_905_2237# m1_2488_2128# m1_1704_1482# li_905_2237# VSUBS sky130_fd_pr__pfet_01v8_X3YSY6
XXM33 VSUBS m1_852_1342# m1_2014_1251# XM33/a_n50_n188# sky130_fd_pr__nfet_01v8_PVEW3M
.ends

.subckt latch_layout m1_1878_998# m1_827_1096# m1_430_1104# m1_822_1732# m1_1595_1096#
+ m1_1097_1325# m1_1878_1968# li_30_2070# m1_1601_1730# m1_724_1961# m1_330_1963#
+ VSUBS
XXM23 VSUBS m1_430_1104# m1_827_1096# m1_1097_1325# sky130_fd_pr__nfet_01v8_PVEW3M
XXM24 VSUBS m1_1595_1096# m1_1097_1325# m1_430_1104# sky130_fd_pr__nfet_01v8_PVEW3M
XXM14 li_30_2070# m1_724_1961# m1_822_1732# li_30_2070# VSUBS sky130_fd_pr__pfet_01v8_X3YSY6
XXM13 li_30_2070# m1_330_1963# m1_430_1104# li_30_2070# VSUBS sky130_fd_pr__pfet_01v8_X3YSY6
XXM15 li_30_2070# m1_1097_1325# m1_430_1104# m1_822_1732# VSUBS sky130_fd_pr__pfet_01v8_X3YSY6
XXM16 li_30_2070# m1_430_1104# m1_1601_1730# m1_1097_1325# VSUBS sky130_fd_pr__pfet_01v8_X3YSY6
XXM17 li_30_2070# m1_1878_1968# li_30_2070# m1_1601_1730# VSUBS sky130_fd_pr__pfet_01v8_X3YSY6
XXM19 VSUBS VSUBS m1_1595_1096# m1_1878_998# sky130_fd_pr__nfet_01v8_PVEW3M
Xsky130_fd_pr__pfet_01v8_X3YSY6_0 li_30_2070# m1_1878_998# li_30_2070# m1_1097_1325#
+ VSUBS sky130_fd_pr__pfet_01v8_X3YSY6
XXM20 VSUBS VSUBS m1_1097_1325# m1_1878_1968# sky130_fd_pr__nfet_01v8_PVEW3M
XXM21 VSUBS m1_430_1104# VSUBS m1_724_1961# sky130_fd_pr__nfet_01v8_PVEW3M
XXM22 VSUBS m1_827_1096# VSUBS m1_330_1963# sky130_fd_pr__nfet_01v8_PVEW3M
.ends

.subckt comparator_full_compact Vdd clk Vc- V+ V- Vc+ Q Q1 m1_2098_364# latch_layout_0/m1_827_1096#
+ vo1- latch_layout_0/m1_1595_1096# latch_layout_0/m1_822_1732# latch_layout_0/m1_1601_1730#
+ comparator_layout_0/m1_852_1342# m1_950_364# vo- vo1+ gnd vo+
Xinverter_0 vo- vo1- Vdd gnd inverter
Xinverter_1 vo+ vo1+ Vdd gnd inverter
Xcomparator_layout_0 vo- vo+ clk Vdd m1_2098_364# V- Vc- m1_950_364# comparator_layout_0/m1_852_1342#
+ gnd Vc+ V+ comparator_layout
Xlatch_layout_0 vo+ latch_layout_0/m1_827_1096# Q latch_layout_0/m1_822_1732# latch_layout_0/m1_1595_1096#
+ Q1 vo1- Vdd latch_layout_0/m1_1601_1730# vo1+ vo- gnd latch_layout
.ends

.subckt sky130_fd_pr__pfet_01v8_lvt_T5G9WD a_n108_n64# w_n144_n164# a_50_n64# a_n50_n161#
+ VSUBS
X0 a_50_n64# a_n50_n161# a_n108_n64# w_n144_n164# sky130_fd_pr__pfet_01v8_lvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
.ends

.subckt sky130_fd_pr__pfet_01v8_lvt_46RJ2R w_n494_n164# a_400_n64# a_n400_n161# a_n458_n64#
+ VSUBS
X0 a_400_n64# a_n400_n161# a_n458_n64# w_n494_n164# sky130_fd_pr__pfet_01v8_lvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=4
.ends

.subckt reference Vdd gnd vo1 vo2 VSUBS
Xsky130_fd_pr__pfet_01v8_lvt_T5G9WD_0 vo1 vo2 vo2 vo1 VSUBS sky130_fd_pr__pfet_01v8_lvt_T5G9WD
Xsky130_fd_pr__pfet_01v8_lvt_46RJ2R_0 Vdd vo2 vo2 Vdd VSUBS sky130_fd_pr__pfet_01v8_lvt_46RJ2R
Xsky130_fd_pr__pfet_01v8_lvt_46RJ2R_1 vo1 vo1 gnd gnd VSUBS sky130_fd_pr__pfet_01v8_lvt_46RJ2R
.ends

.subckt sky130_fd_sc_hd__xnor2_4 A B VGND VNB VPB VPWR Y a_38_47# a_902_47# a_820_297#
+ a_38_297#
X0 VGND A a_902_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1 Y a_38_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2 a_38_297# B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3 a_820_297# B Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4 VPWR a_38_297# Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=2.56 w=1 l=0.15
X5 VGND A a_902_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X6 VGND B a_902_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X7 VGND B a_902_47# VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X8 Y B a_820_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X9 a_38_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X10 a_38_297# B a_38_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X11 VGND A a_38_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X12 a_902_47# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X13 a_820_297# B Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X14 a_902_47# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X15 VPWR A a_38_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X16 Y a_38_297# a_902_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X17 Y a_38_297# a_902_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X18 a_38_47# B a_38_297# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X19 a_38_47# B a_38_297# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X20 a_38_297# B a_38_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.182 ps=1.86 w=0.65 l=0.15
X21 a_38_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X22 VPWR B a_38_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=2.56 w=1 l=0.15
X23 a_38_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X24 a_902_47# a_38_297# Y VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X25 a_902_47# a_38_297# Y VNB sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.0878 ps=0.92 w=0.65 l=0.15
X26 Y B a_820_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X27 a_38_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X28 a_820_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X29 VPWR A a_38_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X30 VGND A a_38_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X31 VPWR A a_820_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X32 a_902_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X33 a_820_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X34 Y a_38_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.135 ps=1.27 w=1 l=0.15
X35 a_902_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X36 a_38_297# B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X37 VPWR A a_820_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X38 VPWR a_38_297# Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X39 VPWR B a_38_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
.ends

.subckt xnor B A gnd Y sky130_fd_sc_hd__xnor2_4_0/a_38_297# sky130_fd_sc_hd__xnor2_4_0/a_38_47#
+ sky130_fd_sc_hd__xnor2_4_0/a_820_297# sky130_fd_sc_hd__xnor2_4_0/VPB Vdd sky130_fd_sc_hd__xnor2_4_0/a_902_47#
+ VSUBS
Xsky130_fd_sc_hd__xnor2_4_0 A B gnd VSUBS sky130_fd_sc_hd__xnor2_4_0/VPB Vdd Y sky130_fd_sc_hd__xnor2_4_0/a_38_47#
+ sky130_fd_sc_hd__xnor2_4_0/a_902_47# sky130_fd_sc_hd__xnor2_4_0/a_820_297# sky130_fd_sc_hd__xnor2_4_0/a_38_297#
+ sky130_fd_sc_hd__xnor2_4
.ends


Xsky130_fd_pr__nfet_01v8_GWFSUW_1 Vdd gnd Vdd gnd gnd Vdd gnd gnd Vdd Vdd gnd Vdd
+ Vdd gnd Vdd gnd gnd gnd sky130_fd_pr__nfet_01v8_GWFSUW
Xcomparator_full_compact_1 Vdd clk Vc+ V+ V- Vc- q comparator_full_compact_1/Q1 comparator_full_compact_1/m1_2098_364#
+ comparator_full_compact_1/latch_layout_0/m1_827_1096# comparator_full_compact_1/vo1-
+ comparator_full_compact_1/latch_layout_0/m1_1595_1096# comparator_full_compact_1/latch_layout_0/m1_822_1732#
+ comparator_full_compact_1/latch_layout_0/m1_1601_1730# comparator_full_compact_1/comparator_layout_0/m1_852_1342#
+ comparator_full_compact_1/m1_950_364# comparator_full_compact_1/vo- comparator_full_compact_1/vo1+
+ gnd comparator_full_compact_1/vo+ comparator_full_compact
Xsky130_fd_pr__nfet_01v8_GWFSUW_2 Vdd gnd Vdd gnd gnd Vdd gnd gnd Vdd Vdd gnd Vdd
+ Vdd gnd Vdd gnd gnd gnd sky130_fd_pr__nfet_01v8_GWFSUW
Xsky130_fd_pr__nfet_01v8_GWFSUW_4 Vdd gnd Vdd gnd gnd Vdd gnd gnd Vdd Vdd gnd Vdd
+ Vdd gnd Vdd gnd gnd gnd sky130_fd_pr__nfet_01v8_GWFSUW
Xsky130_fd_pr__nfet_01v8_GWFSUW_3 Vdd gnd Vdd gnd gnd Vdd gnd gnd Vdd Vdd gnd Vdd
+ Vdd gnd Vdd gnd gnd gnd sky130_fd_pr__nfet_01v8_GWFSUW
Xsky130_fd_pr__nfet_01v8_GWFSUW_5 Vdd gnd Vdd gnd gnd Vdd gnd gnd Vdd Vdd gnd Vdd
+ Vdd gnd Vdd gnd gnd gnd sky130_fd_pr__nfet_01v8_GWFSUW
Xreference_0 Vdd gnd Vc- Vc+ gnd reference
Xxnor_0 q2 q gnd enable xnor_0/sky130_fd_sc_hd__xnor2_4_0/a_38_297# xnor_0/sky130_fd_sc_hd__xnor2_4_0/a_38_47#
+ xnor_0/sky130_fd_sc_hd__xnor2_4_0/a_820_297# xnor_0/sky130_fd_sc_hd__xnor2_4_0/VPB
+ Vdd xnor_0/sky130_fd_sc_hd__xnor2_4_0/a_902_47# gnd xnor
Xcomparator_full_compact_0 Vdd clk Vc- V+ V- Vc+ q2 comparator_full_compact_0/Q1 comparator_full_compact_0/m1_2098_364#
+ comparator_full_compact_0/latch_layout_0/m1_827_1096# comparator_full_compact_0/vo1-
+ comparator_full_compact_0/latch_layout_0/m1_1595_1096# comparator_full_compact_0/latch_layout_0/m1_822_1732#
+ comparator_full_compact_0/latch_layout_0/m1_1601_1730# comparator_full_compact_0/comparator_layout_0/m1_852_1342#
+ comparator_full_compact_0/m1_950_364# comparator_full_compact_0/vo- comparator_full_compact_0/vo1+
+ gnd comparator_full_compact_0/vo+ comparator_full_compact
Xsky130_fd_pr__nfet_01v8_GWFSUW_0 Vdd gnd Vdd gnd gnd Vdd gnd gnd Vdd Vdd gnd Vdd
+ Vdd gnd Vdd gnd gnd gnd sky130_fd_pr__nfet_01v8_GWFSUW


