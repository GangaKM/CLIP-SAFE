* SPICE3 file created from cp1_buffer_5stage.ext - technology: sky130A

X0 cp1_buffer1_0/buffer_digital_0/a_116_148# cp1_buffer1_0/m1_7815_199# cp1_buffer1_2/charge_pump1_0/vdd cp1_buffer1_2/charge_pump1_0/vdd sky130_fd_pr__pfet_01v8 ad=0.365 pd=3.1 as=0.365 ps=3.1 w=1.26 l=0.15
X1 cp1_buffer1_0/charge_pump1_0/clk_in cp1_buffer1_0/buffer_digital_0/a_116_148# cp1_buffer1_2/charge_pump1_0/vdd cp1_buffer1_2/charge_pump1_0/vdd sky130_fd_pr__pfet_01v8 ad=0.365 pd=3.1 as=1.77k ps=15.1k w=1.26 l=0.15
X2 cp1_buffer1_0/buffer_digital_0/a_116_148# cp1_buffer1_0/m1_7815_199# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X3 cp1_buffer1_0/charge_pump1_0/clk_in cp1_buffer1_0/buffer_digital_0/a_116_148# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=887 ps=9.65k w=0.42 l=0.15
X4 cp1_buffer1_0/buffer_digital_1/a_116_148# cp1_buffer1_0/m2_6586_52# cp1_buffer1_2/charge_pump1_0/vdd cp1_buffer1_2/charge_pump1_0/vdd sky130_fd_pr__pfet_01v8 ad=0.365 pd=3.1 as=0 ps=0 w=1.26 l=0.15
X5 cp1_buffer1_0/m1_7815_199# cp1_buffer1_0/buffer_digital_1/a_116_148# cp1_buffer1_2/charge_pump1_0/vdd cp1_buffer1_2/charge_pump1_0/vdd sky130_fd_pr__pfet_01v8 ad=0.365 pd=3.1 as=0 ps=0 w=1.26 l=0.15
X6 cp1_buffer1_0/buffer_digital_1/a_116_148# cp1_buffer1_0/m2_6586_52# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0 ps=0 w=0.42 l=0.15
X7 cp1_buffer1_0/m1_7815_199# cp1_buffer1_0/buffer_digital_1/a_116_148# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0 ps=0 w=0.42 l=0.15
X8 cp1_buffer1_1/buffer_digital_0/a_116_148# cp1_buffer1_1/m1_7815_199# cp1_buffer1_2/charge_pump1_0/vdd cp1_buffer1_2/charge_pump1_0/vdd sky130_fd_pr__pfet_01v8 ad=0.365 pd=3.1 as=0 ps=0 w=1.26 l=0.15
X9 cp1_buffer1_1/charge_pump1_0/clk_in cp1_buffer1_1/buffer_digital_0/a_116_148# cp1_buffer1_2/charge_pump1_0/vdd cp1_buffer1_2/charge_pump1_0/vdd sky130_fd_pr__pfet_01v8 ad=0.365 pd=3.1 as=0 ps=0 w=1.26 l=0.15
X10 cp1_buffer1_1/buffer_digital_0/a_116_148# cp1_buffer1_1/m1_7815_199# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0 ps=0 w=0.42 l=0.15
X11 cp1_buffer1_1/charge_pump1_0/clk_in cp1_buffer1_1/buffer_digital_0/a_116_148# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0 ps=0 w=0.42 l=0.15
X12 cp1_buffer1_1/buffer_digital_1/a_116_148# cp1_buffer1_reverse_0/charge_pump1_reverse_0/clock_1/clk_in cp1_buffer1_2/charge_pump1_0/vdd cp1_buffer1_2/charge_pump1_0/vdd sky130_fd_pr__pfet_01v8 ad=0.365 pd=3.1 as=0 ps=0 w=1.26 l=0.15
X13 cp1_buffer1_1/m1_7815_199# cp1_buffer1_1/buffer_digital_1/a_116_148# cp1_buffer1_2/charge_pump1_0/vdd cp1_buffer1_2/charge_pump1_0/vdd sky130_fd_pr__pfet_01v8 ad=0.365 pd=3.1 as=0 ps=0 w=1.26 l=0.15
X14 cp1_buffer1_1/buffer_digital_1/a_116_148# cp1_buffer1_reverse_0/charge_pump1_reverse_0/clock_1/clk_in VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0 ps=0 w=0.42 l=0.15
X15 cp1_buffer1_1/m1_7815_199# cp1_buffer1_1/buffer_digital_1/a_116_148# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0 ps=0 w=0.42 l=0.15
X16 cp1_buffer1_2/buffer_digital_0/a_116_148# cp1_buffer1_2/m1_7815_199# cp1_buffer1_2/charge_pump1_0/vdd cp1_buffer1_2/charge_pump1_0/vdd sky130_fd_pr__pfet_01v8 ad=0.365 pd=3.1 as=0 ps=0 w=1.26 l=0.15
X17 cp1_buffer1_2/charge_pump1_0/clk_in cp1_buffer1_2/buffer_digital_0/a_116_148# cp1_buffer1_2/charge_pump1_0/vdd cp1_buffer1_2/charge_pump1_0/vdd sky130_fd_pr__pfet_01v8 ad=0.365 pd=3.1 as=0 ps=0 w=1.26 l=0.15
X18 cp1_buffer1_2/buffer_digital_0/a_116_148# cp1_buffer1_2/m1_7815_199# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0 ps=0 w=0.42 l=0.15
X19 cp1_buffer1_2/charge_pump1_0/clk_in cp1_buffer1_2/buffer_digital_0/a_116_148# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0 ps=0 w=0.42 l=0.15
X20 cp1_buffer1_2/buffer_digital_1/a_116_148# cp1_buffer1_reverse_1/charge_pump1_reverse_0/clock_1/clk_in cp1_buffer1_2/charge_pump1_0/vdd cp1_buffer1_2/charge_pump1_0/vdd sky130_fd_pr__pfet_01v8 ad=0.365 pd=3.1 as=0 ps=0 w=1.26 l=0.15
X21 cp1_buffer1_2/m1_7815_199# cp1_buffer1_2/buffer_digital_1/a_116_148# cp1_buffer1_2/charge_pump1_0/vdd cp1_buffer1_2/charge_pump1_0/vdd sky130_fd_pr__pfet_01v8 ad=0.365 pd=3.1 as=0 ps=0 w=1.26 l=0.15
X22 cp1_buffer1_2/buffer_digital_1/a_116_148# cp1_buffer1_reverse_1/charge_pump1_reverse_0/clock_1/clk_in VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0 ps=0 w=0.42 l=0.15
X23 cp1_buffer1_2/m1_7815_199# cp1_buffer1_2/buffer_digital_1/a_116_148# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0 ps=0 w=0.42 l=0.15
X24 cp1_buffer1_reverse_0/buffer_digital_0/a_116_148# cp1_buffer1_reverse_0/m1_7815_199# cp1_buffer1_2/charge_pump1_0/vdd cp1_buffer1_2/charge_pump1_0/vdd sky130_fd_pr__pfet_01v8 ad=0.365 pd=3.1 as=0 ps=0 w=1.26 l=0.15
X25 cp1_buffer1_reverse_0/charge_pump1_reverse_0/clock_1/clk_in cp1_buffer1_reverse_0/buffer_digital_0/a_116_148# cp1_buffer1_2/charge_pump1_0/vdd cp1_buffer1_2/charge_pump1_0/vdd sky130_fd_pr__pfet_01v8 ad=0.365 pd=3.1 as=0 ps=0 w=1.26 l=0.15
X26 cp1_buffer1_reverse_0/buffer_digital_0/a_116_148# cp1_buffer1_reverse_0/m1_7815_199# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0 ps=0 w=0.42 l=0.15
X27 cp1_buffer1_reverse_0/charge_pump1_reverse_0/clock_1/clk_in cp1_buffer1_reverse_0/buffer_digital_0/a_116_148# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0 ps=0 w=0.42 l=0.15
X28 cp1_buffer1_reverse_0/buffer_digital_1/a_116_148# cp1_buffer1_0/charge_pump1_0/clk_in cp1_buffer1_2/charge_pump1_0/vdd cp1_buffer1_2/charge_pump1_0/vdd sky130_fd_pr__pfet_01v8 ad=0.365 pd=3.1 as=0 ps=0 w=1.26 l=0.15
X29 cp1_buffer1_reverse_0/m1_7815_199# cp1_buffer1_reverse_0/buffer_digital_1/a_116_148# cp1_buffer1_2/charge_pump1_0/vdd cp1_buffer1_2/charge_pump1_0/vdd sky130_fd_pr__pfet_01v8 ad=0.365 pd=3.1 as=0 ps=0 w=1.26 l=0.15
X30 cp1_buffer1_reverse_0/buffer_digital_1/a_116_148# cp1_buffer1_0/charge_pump1_0/clk_in VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0 ps=0 w=0.42 l=0.15
X31 cp1_buffer1_reverse_0/m1_7815_199# cp1_buffer1_reverse_0/buffer_digital_1/a_116_148# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0 ps=0 w=0.42 l=0.15
X32 cp1_buffer1_reverse_1/buffer_digital_0/a_116_148# cp1_buffer1_reverse_1/m1_7815_199# cp1_buffer1_2/charge_pump1_0/vdd cp1_buffer1_2/charge_pump1_0/vdd sky130_fd_pr__pfet_01v8 ad=0.365 pd=3.1 as=0 ps=0 w=1.26 l=0.15
X33 cp1_buffer1_reverse_1/charge_pump1_reverse_0/clock_1/clk_in cp1_buffer1_reverse_1/buffer_digital_0/a_116_148# cp1_buffer1_2/charge_pump1_0/vdd cp1_buffer1_2/charge_pump1_0/vdd sky130_fd_pr__pfet_01v8 ad=0.365 pd=3.1 as=0 ps=0 w=1.26 l=0.15
X34 cp1_buffer1_reverse_1/buffer_digital_0/a_116_148# cp1_buffer1_reverse_1/m1_7815_199# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0 ps=0 w=0.42 l=0.15
X35 cp1_buffer1_reverse_1/charge_pump1_reverse_0/clock_1/clk_in cp1_buffer1_reverse_1/buffer_digital_0/a_116_148# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0 ps=0 w=0.42 l=0.15
X36 cp1_buffer1_reverse_1/buffer_digital_1/a_116_148# cp1_buffer1_1/charge_pump1_0/clk_in cp1_buffer1_2/charge_pump1_0/vdd cp1_buffer1_2/charge_pump1_0/vdd sky130_fd_pr__pfet_01v8 ad=0.365 pd=3.1 as=0 ps=0 w=1.26 l=0.15
X37 cp1_buffer1_reverse_1/m1_7815_199# cp1_buffer1_reverse_1/buffer_digital_1/a_116_148# cp1_buffer1_2/charge_pump1_0/vdd cp1_buffer1_2/charge_pump1_0/vdd sky130_fd_pr__pfet_01v8 ad=0.365 pd=3.1 as=0 ps=0 w=1.26 l=0.15
X38 cp1_buffer1_reverse_1/buffer_digital_1/a_116_148# cp1_buffer1_1/charge_pump1_0/clk_in VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0 ps=0 w=0.42 l=0.15
X39 cp1_buffer1_reverse_1/m1_7815_199# cp1_buffer1_reverse_1/buffer_digital_1/a_116_148# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0 ps=0 w=0.42 l=0.15
C0 cp1_buffer1_reverse_1/charge_pump1_reverse_0/capacitors_1_7/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# VSUBS 6.15f
C1 cp1_buffer1_2/charge_pump1_0/clkb cp1_buffer1_2/charge_pump1_0/clock_0/a_2432_n962# 2.67f
C2 cp1_buffer1_reverse_1/charge_pump1_reverse_0/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# cp1_buffer1_2/charge_pump1_0/vdd 3.48f
C3 cp1_buffer1_2/charge_pump1_0/in2 cp1_buffer1_reverse_0/charge_pump1_reverse_0/capacitors_1_10/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 2.94f
C4 VSUBS cp1_buffer1_2/charge_pump1_0/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 6.15f
C5 cp1_buffer1_reverse_1/charge_pump1_reverse_0/capacitors_1_7/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# cp1_buffer1_2/charge_pump1_0/vdd 3.49f
C6 VSUBS cp1_buffer1_2/charge_pump1_0/capacitors_1_9/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 6.15f
C7 cp1_buffer1_2/charge_pump1_0/in2 cp1_buffer1_2/charge_pump1_0/capacitors_1_2/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 2.94f
C8 cp1_buffer1_2/charge_pump1_0/vdd cp1_buffer1_1/charge_pump1_0/capacitor_8_1/capacitor_7_0/buffer_and_gate_0/m1_5444_838# 8.43f
C9 cp1_buffer1_0/charge_pump1_0/capacitors_1_5/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# cp1_buffer1_2/charge_pump1_0/vdd 3.48f
C10 cp1_buffer1_reverse_0/charge_pump1_reverse_0/capacitors_1_4/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/m1_5444_838# cp1_buffer1_2/charge_pump1_0/vdd 8.43f
C11 cp1_buffer1_reverse_0/charge_pump1_reverse_0/capacitors_1_2/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/m1_5444_838# cp1_buffer1_2/charge_pump1_0/vdd 8.44f
C12 cp1_buffer1_1/charge_pump1_0/capacitors_1_12/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/m1_5444_838# VSUBS 4.07f
C13 cp1_buffer1_2/charge_pump1_0/capacitors_1_6/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# cp1_buffer1_2/charge_pump1_0/capacitors_1_6/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/m1_5444_838# 2.1f
C14 cp1_buffer1_0/charge_pump1_0/capacitors_1_2/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# cp1_buffer1_2/charge_pump1_0/vdd 13.3f
C15 cp1_buffer1_0/charge_pump1_0/capacitors_1_12/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# cp1_buffer1_2/charge_pump1_0/vdd 3.48f
C16 cp1_buffer1_reverse_1/charge_pump1_reverse_0/clock_1/clk cp1_buffer1_reverse_1/charge_pump1_reverse_0/capacitors_1_1/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 2.18f
C17 cp1_buffer1_reverse_1/charge_pump1_reverse_0/capacitors_1_13/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# cp1_buffer1_2/charge_pump1_0/vdd 13.3f
C18 cp1_buffer1_1/charge_pump1_0/capacitors_1_11/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# cp1_buffer1_2/charge_pump1_0/vdd 3.49f
C19 cp1_buffer1_0/charge_pump1_0/capacitors_1_10/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# cp1_buffer1_2/charge_pump1_0/vdd 13.3f
C20 cp1_buffer1_reverse_0/charge_pump1_reverse_0/capacitors_1_4/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# VSUBS 6.15f
C21 cp1_buffer1_1/charge_pump1_0/capacitor_8_1/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# cp1_buffer1_1/charge_pump1_0/capacitor_8_1/capacitor_7_0/buffer_and_gate_0/m1_5444_838# 2.1f
C22 cp1_buffer1_reverse_0/charge_pump1_reverse_0/capacitors_1_2/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# VSUBS 6.15f
C23 cp1_buffer1_2/charge_pump1_0/capacitors_1_1/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# cp1_buffer1_2/charge_pump1_0/vdd 13.1f
C24 cp1_buffer1_0/charge_pump1_0/capacitors_1_8/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/m1_5444_838# cp1_buffer1_2/charge_pump1_0/vdd 8.44f
C25 cp1_buffer1_reverse_0/charge_pump1_reverse_0/capacitors_1_4/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# cp1_buffer1_2/charge_pump1_0/vdd 3.48f
C26 cp1_buffer1_reverse_0/charge_pump1_reverse_0/capacitors_1_2/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# cp1_buffer1_2/charge_pump1_0/vdd 3.49f
C27 VSUBS cp1_buffer1_1/charge_pump1_0/capacitors_1_1/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/m1_5444_838# 4f
C28 cp1_buffer1_reverse_0/charge_pump1_reverse_0/input2 cp1_buffer1_reverse_0/charge_pump1_reverse_0/clock_1/clk 8.93f
C29 cp1_buffer1_2/charge_pump1_0/in2 VSUBS 7.32f
C30 cp1_buffer1_2/charge_pump1_0/capacitors_1_11/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 cp1_buffer1_2/charge_pump1_0/in6 2.94f
C31 cp1_buffer1_1/charge_pump1_0/capacitors_1_11/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/m1_5444_838# VSUBS 4.08f
C32 VSUBS cp1_buffer1_1/charge_pump1_0/capacitors_1_9/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 6.15f
C33 cp1_buffer1_reverse_1/charge_pump1_reverse_0/capacitors_1_4/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 cp1_buffer1_2/charge_pump1_0/in7 2.94f
C34 cp1_buffer1_reverse_0/charge_pump1_reverse_0/capacitor_8_1/capacitor_7_0/buffer_and_gate_0/m1_5444_838# cp1_buffer1_reverse_0/charge_pump1_reverse_0/capacitor_8_1/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 2.1f
C35 cp1_buffer1_reverse_1/charge_pump1_reverse_0/capacitors_1_1/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/m1_5444_838# cp1_buffer1_2/charge_pump1_0/vdd 8.43f
C36 cp1_buffer1_2/charge_pump1_0/capacitor_8_1/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# cp1_buffer1_2/charge_pump1_0/vdd 13.3f
C37 cp1_buffer1_0/charge_pump1_0/capacitor_8_1/capacitor_7_0/buffer_and_gate_0/m1_5444_838# VSUBS 4.07f
C38 cp1_buffer1_reverse_1/charge_pump1_reverse_0/capacitors_1_12/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/m1_5444_838# VSUBS 4.07f
C39 cp1_buffer1_1/charge_pump1_0/capacitors_1_10/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/m1_5444_838# VSUBS 4.07f
C40 cp1_buffer1_2/charge_pump1_0/clkb cp1_buffer1_2/charge_pump1_0/g2 8.12f
C41 cp1_buffer1_reverse_1/charge_pump1_reverse_0/capacitors_1_1/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# VSUBS 6.05f
C42 cp1_buffer1_reverse_1/charge_pump1_reverse_0/clock_1/clk cp1_buffer1_reverse_1/charge_pump1_reverse_0/capacitors_1_11/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 2.16f
C43 cp1_buffer1_reverse_0/charge_pump1_reverse_0/clock_1/a_2020_n482# cp1_buffer1_2/charge_pump1_0/vdd 2.66f
C44 cp1_buffer1_0/charge_pump1_0/clk cp1_buffer1_0/charge_pump1_0/capacitors_1_7/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 2.17f
C45 cp1_buffer1_reverse_0/charge_pump1_reverse_0/capacitors_1_1/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# cp1_buffer1_2/charge_pump1_0/vdd 13.1f
C46 cp1_buffer1_reverse_0/charge_pump1_reverse_0/capacitor_8_1/capacitor_7_0/buffer_and_gate_0/m1_5444_838# cp1_buffer1_2/charge_pump1_0/vdd 8.43f
C47 cp1_buffer1_2/charge_pump1_0/in1 cp1_buffer1_2/charge_pump1_0/vdd 14f
C48 cp1_buffer1_reverse_1/charge_pump1_reverse_0/capacitors_1_1/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# cp1_buffer1_2/charge_pump1_0/vdd 3.45f
C49 cp1_buffer1_2/charge_pump1_0/capacitors_1_7/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/m1_5444_838# cp1_buffer1_2/charge_pump1_0/capacitors_1_7/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 2.1f
C50 cp1_buffer1_0/charge_pump1_0/capacitors_1_1/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/m1_5444_838# cp1_buffer1_2/charge_pump1_0/vdd 8.43f
C51 cp1_buffer1_reverse_1/charge_pump1_reverse_0/capacitors_1_9/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# cp1_buffer1_2/charge_pump1_0/vdd 13.3f
C52 cp1_buffer1_reverse_0/charge_pump1_reverse_0/capacitors_1_6/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# cp1_buffer1_2/charge_pump1_0/vdd 13.3f
C53 cp1_buffer1_2/charge_pump1_0/capacitors_1_10/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/m1_5444_838# VSUBS 4.07f
C54 cp1_buffer1_2/charge_pump1_0/in4 cp1_buffer1_2/charge_pump1_0/capacitors_1_6/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 2.94f
C55 cp1_buffer1_2/charge_pump1_0/capacitors_1_0/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# cp1_buffer1_2/charge_pump1_0/vdd 3.45f
C56 cp1_buffer1_reverse_0/charge_pump1_reverse_0/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# cp1_buffer1_2/charge_pump1_0/vdd 13.3f
C57 cp1_buffer1_0/charge_pump1_0/capacitors_1_7/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/m1_5444_838# cp1_buffer1_0/charge_pump1_0/capacitors_1_7/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 2.1f
C58 cp1_buffer1_reverse_1/charge_pump1_reverse_0/capacitors_1_11/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/m1_5444_838# cp1_buffer1_2/charge_pump1_0/vdd 8.44f
C59 cp1_buffer1_2/charge_pump1_0/vdd cp1_buffer1_1/charge_pump1_0/clock_0/a_3246_118# 7.35f
C60 cp1_buffer1_reverse_0/charge_pump1_reverse_0/capacitors_1_3/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/m1_5444_838# VSUBS 4.07f
C61 cp1_buffer1_2/charge_pump1_0/vdd cp1_buffer1_1/charge_pump1_0/capacitors_1_5/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 13.3f
C62 VSUBS cp1_buffer1_1/charge_pump1_0/capacitors_1_7/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 6.15f
C63 cp1_buffer1_0/charge_pump1_0/g1 cp1_buffer1_0/charge_pump1_0/clk 8.15f
C64 cp1_buffer1_1/charge_pump1_0/clkb cp1_buffer1_1/charge_pump1_0/input2 8.93f
C65 cp1_buffer1_reverse_1/charge_pump1_reverse_0/capacitors_1_11/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# VSUBS 6.15f
C66 cp1_buffer1_2/charge_pump1_0/input2 cp1_buffer1_2/charge_pump1_0/input1 3.33f
C67 cp1_buffer1_2/charge_pump1_0/in8 cp1_buffer1_2/charge_pump1_0/vdd 13.6f
C68 cp1_buffer1_reverse_1/charge_pump1_reverse_0/capacitors_1_11/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# cp1_buffer1_2/charge_pump1_0/vdd 3.49f
C69 cp1_buffer1_2/charge_pump1_0/capacitors_1_5/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# cp1_buffer1_2/charge_pump1_0/clkb 2.16f
C70 cp1_buffer1_2/charge_pump1_0/in1 cp1_buffer1_0/charge_pump1_0/capacitors_1_0/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 2.94f
C71 VSUBS cp1_buffer1_2/charge_pump1_0/capacitors_1_7/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 6.15f
C72 VSUBS cp1_buffer1_1/charge_pump1_0/capacitors_1_2/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 6.15f
C73 cp1_buffer1_reverse_1/charge_pump1_reverse_0/capacitors_1_3/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# cp1_buffer1_reverse_1/charge_pump1_reverse_0/capacitors_1_3/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/m1_5444_838# 2.1f
C74 cp1_buffer1_reverse_0/charge_pump1_reverse_0/clock_1/clkb cp1_buffer1_2/charge_pump1_0/vdd 83.4f
C75 cp1_buffer1_1/charge_pump1_0/capacitors_1_3/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# VSUBS 6.15f
C76 cp1_buffer1_reverse_1/charge_pump1_reverse_0/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# cp1_buffer1_reverse_1/charge_pump1_reverse_0/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/m1_5444_838# 2.1f
C77 cp1_buffer1_2/charge_pump1_0/capacitors_1_4/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# cp1_buffer1_2/charge_pump1_0/capacitors_1_4/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/m1_5444_838# 2.1f
C78 cp1_buffer1_1/charge_pump1_0/capacitors_1_0/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# cp1_buffer1_2/charge_pump1_0/vdd 13.1f
C79 cp1_buffer1_0/charge_pump1_0/m1_4341_n519# cp1_buffer1_0/charge_pump1_0/clk 9.42f
C80 cp1_buffer1_reverse_1/charge_pump1_reverse_0/clock_1/a_2020_n482# cp1_buffer1_2/charge_pump1_0/vdd 2.66f
C81 cp1_buffer1_reverse_1/charge_pump1_reverse_0/capacitors_1_5/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 cp1_buffer1_2/charge_pump1_0/in6 2.94f
C82 cp1_buffer1_1/charge_pump1_0/m1_12659_300# cp1_buffer1_1/charge_pump1_0/clkb 9.47f
C83 cp1_buffer1_2/charge_pump1_0/capacitors_1_9/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/m1_5444_838# VSUBS 4.07f
C84 cp1_buffer1_reverse_1/charge_pump1_reverse_0/capacitors_1_12/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# cp1_buffer1_reverse_1/charge_pump1_reverse_0/capacitors_1_12/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/m1_5444_838# 2.1f
C85 cp1_buffer1_2/charge_pump1_0/capacitors_1_5/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/m1_5444_838# VSUBS 4.07f
C86 cp1_buffer1_2/charge_pump1_0/vdd cp1_buffer1_1/charge_pump1_0/capacitors_1_11/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 13.3f
C87 cp1_buffer1_0/charge_pump1_0/capacitors_1_8/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 cp1_buffer1_2/charge_pump1_0/in6 2.94f
C88 cp1_buffer1_reverse_1/charge_pump1_reverse_0/capacitors_1_2/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/m1_5444_838# VSUBS 4.07f
C89 cp1_buffer1_1/charge_pump1_0/capacitors_1_13/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# cp1_buffer1_2/charge_pump1_0/vdd 3.48f
C90 cp1_buffer1_reverse_0/charge_pump1_reverse_0/capacitors_1_5/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/m1_5444_838# cp1_buffer1_2/charge_pump1_0/vdd 8.44f
C91 cp1_buffer1_2/charge_pump1_0/capacitors_1_8/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/m1_5444_838# VSUBS 4.07f
C92 cp1_buffer1_1/charge_pump1_0/clkb cp1_buffer1_1/charge_pump1_0/g2 8.12f
C93 cp1_buffer1_2/charge_pump1_0/vdd cp1_buffer1_0/charge_pump1_0/capacitors_1_7/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 13.3f
C94 cp1_buffer1_reverse_0/charge_pump1_reverse_0/capacitors_1_5/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# VSUBS 6.15f
C95 cp1_buffer1_reverse_0/charge_pump1_reverse_0/input2 cp1_buffer1_2/charge_pump1_0/vdd 28f
C96 cp1_buffer1_reverse_1/charge_pump1_reverse_0/capacitors_1_4/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# cp1_buffer1_2/charge_pump1_0/vdd 13.3f
C97 cp1_buffer1_reverse_1/charge_pump1_reverse_0/input2 cp1_buffer1_reverse_1/charge_pump1_reverse_0/input1 3.33f
C98 cp1_buffer1_reverse_1/charge_pump1_reverse_0/capacitors_1_9/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 cp1_buffer1_2/charge_pump1_0/in2 2.94f
C99 cp1_buffer1_reverse_1/charge_pump1_reverse_0/clock_1/clkb VSUBS 28.4f
C100 cp1_buffer1_reverse_1/charge_pump1_reverse_0/capacitors_1_10/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/m1_5444_838# VSUBS 4.07f
C101 cp1_buffer1_reverse_0/charge_pump1_reverse_0/capacitors_1_5/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# cp1_buffer1_2/charge_pump1_0/vdd 3.48f
C102 cp1_buffer1_1/charge_pump1_0/capacitors_1_13/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/m1_5444_838# VSUBS 4.07f
C103 cp1_buffer1_2/charge_pump1_0/in2 cp1_buffer1_1/charge_pump1_0/capacitors_1_4/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 2.94f
C104 cp1_buffer1_1/charge_pump1_0/capacitors_1_8/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/m1_5444_838# cp1_buffer1_2/charge_pump1_0/vdd 8.44f
C105 cp1_buffer1_reverse_1/charge_pump1_reverse_0/capacitor_8_1/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# cp1_buffer1_2/charge_pump1_0/vdd 13.3f
C106 cp1_buffer1_2/charge_pump1_0/capacitor_8_1/capacitor_7_0/buffer_and_gate_0/m1_5444_838# cp1_buffer1_2/charge_pump1_0/vdd 8.43f
C107 cp1_buffer1_reverse_0/charge_pump1_reverse_0/m1_12659_300# cp1_buffer1_1/charge_pump1_0/vin 2.14f
C108 cp1_buffer1_0/charge_pump1_0/capacitors_1_2/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/m1_5444_838# VSUBS 4.07f
C109 cp1_buffer1_reverse_1/charge_pump1_reverse_0/clock_1/clk cp1_buffer1_reverse_1/charge_pump1_reverse_0/nmos_dnw3_0/clkb 8.35f
C110 cp1_buffer1_1/charge_pump1_0/clk cp1_buffer1_1/charge_pump1_0/clock_0/a_3246_118# 2.71f
C111 cp1_buffer1_2/charge_pump1_0/vdd cp1_buffer1_1/charge_pump1_0/capacitors_1_7/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/m1_5444_838# 8.44f
C112 cp1_buffer1_2/charge_pump1_0/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/m1_5444_838# cp1_buffer1_2/charge_pump1_0/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 2.1f
C113 cp1_buffer1_2/charge_pump1_0/clk_in VSUBS 3.43f
C114 cp1_buffer1_reverse_1/charge_pump1_reverse_0/clock_1/a_3246_118# cp1_buffer1_2/charge_pump1_0/vdd 7.37f
C115 cp1_buffer1_0/charge_pump1_0/capacitors_1_4/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/m1_5444_838# cp1_buffer1_0/charge_pump1_0/capacitors_1_4/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 2.1f
C116 cp1_buffer1_0/charge_pump1_0/capacitors_1_3/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/m1_5444_838# cp1_buffer1_0/charge_pump1_0/capacitors_1_3/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 2.1f
C117 cp1_buffer1_reverse_0/charge_pump1_reverse_0/clock_1/clkb cp1_buffer1_reverse_0/charge_pump1_reverse_0/clock_1/a_2432_n962# 2.69f
C118 cp1_buffer1_1/charge_pump1_0/capacitors_1_10/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# cp1_buffer1_2/charge_pump1_0/vdd 13.3f
C119 cp1_buffer1_0/charge_pump1_0/capacitors_1_11/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/m1_5444_838# cp1_buffer1_2/charge_pump1_0/vdd 8.44f
C120 cp1_buffer1_2/charge_pump1_0/capacitors_1_3/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# cp1_buffer1_2/charge_pump1_0/capacitors_1_3/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/m1_5444_838# 2.1f
C121 cp1_buffer1_2/charge_pump1_0/capacitors_1_2/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# cp1_buffer1_2/charge_pump1_0/vdd 3.49f
C122 cp1_buffer1_2/charge_pump1_0/vdd cp1_buffer1_1/charge_pump1_0/capacitors_1_4/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 13.3f
C123 cp1_buffer1_1/charge_pump1_0/clk_in VSUBS 6.42f
C124 cp1_buffer1_2/charge_pump1_0/vdd cp1_buffer1_2/charge_pump1_0/capacitors_1_3/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/m1_5444_838# 8.44f
C125 cp1_buffer1_reverse_0/charge_pump1_reverse_0/capacitors_1_3/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# cp1_buffer1_reverse_0/charge_pump1_reverse_0/capacitors_1_3/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/m1_5444_838# 2.1f
C126 cp1_buffer1_1/charge_pump1_0/capacitors_1_0/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# cp1_buffer1_1/charge_pump1_0/capacitors_1_0/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/m1_5444_838# 2.1f
C127 cp1_buffer1_2/charge_pump1_0/input1 cp1_buffer1_2/charge_pump1_0/clk 8.87f
C128 cp1_buffer1_2/charge_pump1_0/capacitors_1_13/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# cp1_buffer1_2/charge_pump1_0/vdd 13.3f
C129 cp1_buffer1_reverse_0/charge_pump1_reverse_0/capacitors_1_11/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# cp1_buffer1_reverse_0/charge_pump1_reverse_0/clock_1/clk 2.16f
C130 cp1_buffer1_reverse_0/charge_pump1_reverse_0/capacitors_1_9/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# cp1_buffer1_2/charge_pump1_0/vdd 13.3f
C131 cp1_buffer1_0/charge_pump1_0/capacitors_1_12/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# cp1_buffer1_0/charge_pump1_0/capacitors_1_12/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/m1_5444_838# 2.1f
C132 cp1_buffer1_2/charge_pump1_0/clock_0/a_2402_572# cp1_buffer1_2/charge_pump1_0/vdd 2.67f
C133 cp1_buffer1_1/charge_pump1_0/capacitors_1_2/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/m1_5444_838# VSUBS 4.07f
C134 cp1_buffer1_1/charge_pump1_0/capacitors_1_0/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# cp1_buffer1_1/charge_pump1_0/clk 2.2f
C135 cp1_buffer1_reverse_0/charge_pump1_reverse_0/capacitors_1_7/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# cp1_buffer1_2/charge_pump1_0/vdd 13.3f
C136 cp1_buffer1_0/charge_pump1_0/capacitors_1_4/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/m1_5444_838# cp1_buffer1_2/charge_pump1_0/vdd 8.44f
C137 cp1_buffer1_1/charge_pump1_0/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/m1_5444_838# cp1_buffer1_2/charge_pump1_0/vdd 8.43f
C138 cp1_buffer1_2/charge_pump1_0/input2 cp1_buffer1_2/charge_pump1_0/clkb 8.93f
C139 cp1_buffer1_reverse_0/charge_pump1_reverse_0/clock_1/clkb cp1_buffer1_reverse_0/charge_pump1_reverse_0/input1 8.86f
C140 cp1_buffer1_2/charge_pump1_0/capacitors_1_0/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# cp1_buffer1_2/charge_pump1_0/vdd 13.1f
C141 cp1_buffer1_reverse_1/charge_pump1_reverse_0/capacitors_1_8/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 cp1_buffer1_2/charge_pump1_0/in3 2.94f
C142 cp1_buffer1_0/charge_pump1_0/capacitors_1_0/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# cp1_buffer1_2/charge_pump1_0/vdd 3.45f
C143 cp1_buffer1_reverse_0/charge_pump1_reverse_0/capacitors_1_0/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# cp1_buffer1_reverse_0/charge_pump1_reverse_0/capacitors_1_0/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/m1_5444_838# 2.1f
C144 VSUBS cp1_buffer1_reverse_0/charge_pump1_reverse_0/clock_1/clk 30.9f
C145 cp1_buffer1_2/charge_pump1_0/capacitors_1_11/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# cp1_buffer1_2/charge_pump1_0/vdd 13.3f
C146 cp1_buffer1_reverse_1/charge_pump1_reverse_0/capacitors_1_3/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/m1_5444_838# cp1_buffer1_2/charge_pump1_0/vdd 8.44f
C147 cp1_buffer1_0/charge_pump1_0/capacitors_1_5/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# VSUBS 6.15f
C148 cp1_buffer1_0/charge_pump1_0/capacitors_1_6/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# cp1_buffer1_0/charge_pump1_0/clk 2.17f
C149 cp1_buffer1_reverse_0/charge_pump1_reverse_0/capacitors_1_12/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# cp1_buffer1_reverse_0/charge_pump1_reverse_0/capacitors_1_12/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/m1_5444_838# 2.1f
C150 VSUBS cp1_buffer1_1/charge_pump1_0/capacitors_1_9/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/m1_5444_838# 4.07f
C151 cp1_buffer1_2/charge_pump1_0/capacitors_1_4/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/m1_5444_838# VSUBS 4.07f
C152 cp1_buffer1_2/charge_pump1_0/in1 cp1_buffer1_reverse_0/charge_pump1_reverse_0/capacitor_8_1/capacitor_7_0/buffer_and_gate_0/in1 2.94f
C153 cp1_buffer1_2/charge_pump1_0/capacitors_1_4/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# cp1_buffer1_2/charge_pump1_0/vdd 13.3f
C154 cp1_buffer1_0/charge_pump1_0/clkb VSUBS 27.7f
C155 cp1_buffer1_reverse_1/charge_pump1_reverse_0/capacitors_1_3/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# VSUBS 6.15f
C156 cp1_buffer1_2/charge_pump1_0/vdd cp1_buffer1_2/charge_pump1_0/capacitors_1_5/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# 3.48f
C157 cp1_buffer1_1/charge_pump1_0/capacitors_1_7/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# cp1_buffer1_2/charge_pump1_0/vdd 3.49f
C158 cp1_buffer1_1/charge_pump1_0/clock_0/a_2432_n962# cp1_buffer1_2/charge_pump1_0/vdd 7.04f
C159 cp1_buffer1_reverse_1/charge_pump1_reverse_0/capacitors_1_3/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# cp1_buffer1_2/charge_pump1_0/vdd 3.48f
C160 cp1_buffer1_0/charge_pump1_0/capacitors_1_2/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# cp1_buffer1_2/charge_pump1_0/vdd 3.49f
C161 cp1_buffer1_reverse_0/charge_pump1_reverse_0/capacitors_1_3/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 cp1_buffer1_2/charge_pump1_0/in6 2.94f
C162 cp1_buffer1_2/charge_pump1_0/capacitors_1_9/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 cp1_buffer1_2/charge_pump1_0/in7 2.94f
C163 cp1_buffer1_0/charge_pump1_0/capacitors_1_13/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# VSUBS 6.15f
C164 cp1_buffer1_2/charge_pump1_0/in2 cp1_buffer1_1/charge_pump1_0/capacitors_1_2/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 2.94f
C165 cp1_buffer1_0/charge_pump1_0/clk VSUBS 31.5f
C166 cp1_buffer1_reverse_0/charge_pump1_reverse_0/input2 cp1_buffer1_reverse_0/charge_pump1_reverse_0/input1 3.33f
C167 cp1_buffer1_2/charge_pump1_0/capacitors_1_10/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# VSUBS 6.15f
C168 cp1_buffer1_reverse_1/charge_pump1_reverse_0/capacitors_1_0/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/m1_5444_838# cp1_buffer1_2/charge_pump1_0/vdd 8.43f
C169 cp1_buffer1_2/charge_pump1_0/capacitors_1_8/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# cp1_buffer1_2/charge_pump1_0/clk 2.17f
C170 cp1_buffer1_2/charge_pump1_0/capacitors_1_6/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# cp1_buffer1_2/charge_pump1_0/clk 2.17f
C171 cp1_buffer1_2/charge_pump1_0/m1_4341_n519# cp1_buffer1_2/charge_pump1_0/clk 9.42f
C172 VSUBS cp1_buffer1_0/charge_pump1_0/capacitors_1_7/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/m1_5444_838# 4.07f
C173 cp1_buffer1_0/charge_pump1_0/capacitors_1_10/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# cp1_buffer1_2/charge_pump1_0/vdd 3.48f
C174 cp1_buffer1_reverse_1/charge_pump1_reverse_0/clock_1/clk_in VSUBS 5.72f
C175 cp1_buffer1_reverse_0/charge_pump1_reverse_0/capacitors_1_12/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/m1_5444_838# cp1_buffer1_2/charge_pump1_0/vdd 8.44f
C176 VSUBS cp1_buffer1_1/charge_pump1_0/capacitors_1_13/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 6.15f
C177 cp1_buffer1_reverse_0/charge_pump1_reverse_0/clock_1/a_3246_118# cp1_buffer1_reverse_0/charge_pump1_reverse_0/clock_1/clk 2.73f
C178 cp1_buffer1_1/charge_pump1_0/clock_0/a_2020_n482# cp1_buffer1_2/charge_pump1_0/vdd 2.66f
C179 cp1_buffer1_1/charge_pump1_0/capacitors_1_3/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# cp1_buffer1_2/charge_pump1_0/vdd 3.48f
C180 cp1_buffer1_reverse_1/charge_pump1_reverse_0/capacitors_1_5/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# cp1_buffer1_2/charge_pump1_0/vdd 13.3f
C181 cp1_buffer1_reverse_0/charge_pump1_reverse_0/capacitors_1_12/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# VSUBS 6.15f
C182 cp1_buffer1_reverse_1/charge_pump1_reverse_0/capacitors_1_2/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# cp1_buffer1_reverse_1/charge_pump1_reverse_0/capacitors_1_2/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/m1_5444_838# 2.1f
C183 VSUBS cp1_buffer1_1/charge_pump1_0/capacitors_1_1/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 6.05f
C184 cp1_buffer1_0/charge_pump1_0/clock_0/a_2402_572# cp1_buffer1_2/charge_pump1_0/vdd 2.67f
C185 VSUBS cp1_buffer1_0/charge_pump1_0/capacitor_8_1/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 6.15f
C186 VSUBS cp1_buffer1_2/charge_pump1_0/capacitors_1_1/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/m1_5444_838# 4f
C187 cp1_buffer1_reverse_0/charge_pump1_reverse_0/capacitors_1_12/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# cp1_buffer1_2/charge_pump1_0/vdd 3.48f
C188 cp1_buffer1_0/charge_pump1_0/clkb cp1_buffer1_0/charge_pump1_0/capacitors_1_11/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 2.16f
C189 cp1_buffer1_1/charge_pump1_0/clk cp1_buffer1_1/charge_pump1_0/g1 8.15f
C190 cp1_buffer1_2/charge_pump1_0/capacitors_1_7/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/m1_5444_838# cp1_buffer1_2/charge_pump1_0/vdd 8.44f
C191 cp1_buffer1_0/charge_pump1_0/capacitors_1_13/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/m1_5444_838# VSUBS 4.07f
C192 cp1_buffer1_2/charge_pump1_0/in4 cp1_buffer1_1/charge_pump1_0/capacitors_1_13/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 2.94f
C193 cp1_buffer1_0/charge_pump1_0/clk_in cp1_buffer1_2/charge_pump1_0/vdd 7.32f
C194 VSUBS cp1_buffer1_0/charge_pump1_0/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/m1_5444_838# 4.07f
C195 cp1_buffer1_0/charge_pump1_0/clk cp1_buffer1_0/charge_pump1_0/capacitors_1_9/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 2.17f
C196 cp1_buffer1_reverse_1/charge_pump1_reverse_0/clock_1/clk cp1_buffer1_2/charge_pump1_0/vdd 78.8f
C197 cp1_buffer1_2/charge_pump1_0/capacitors_1_10/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 cp1_buffer1_2/charge_pump1_0/in7 2.94f
C198 cp1_buffer1_0/charge_pump1_0/capacitors_1_4/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# VSUBS 6.15f
C199 cp1_buffer1_1/charge_pump1_0/input1 VSUBS 9.98f
C200 cp1_buffer1_reverse_1/charge_pump1_reverse_0/capacitors_1_2/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# cp1_buffer1_reverse_1/charge_pump1_reverse_0/clock_1/clkb 2.17f
C201 cp1_buffer1_reverse_0/charge_pump1_reverse_0/capacitors_1_6/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# cp1_buffer1_reverse_0/charge_pump1_reverse_0/clock_1/clkb 2.17f
C202 cp1_buffer1_0/charge_pump1_0/capacitors_1_6/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# cp1_buffer1_2/charge_pump1_0/vdd 13.3f
C203 cp1_buffer1_reverse_0/charge_pump1_reverse_0/capacitors_1_11/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# cp1_buffer1_2/charge_pump1_0/vdd 13.3f
C204 cp1_buffer1_1/charge_pump1_0/capacitors_1_6/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/m1_5444_838# cp1_buffer1_2/charge_pump1_0/vdd 8.43f
C205 cp1_buffer1_2/charge_pump1_0/capacitors_1_8/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# cp1_buffer1_2/charge_pump1_0/vdd 3.49f
C206 cp1_buffer1_reverse_0/charge_pump1_reverse_0/clock_1/clkb cp1_buffer1_reverse_0/charge_pump1_reverse_0/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 2.17f
C207 cp1_buffer1_reverse_1/charge_pump1_reverse_0/capacitors_1_6/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/m1_5444_838# VSUBS 4.07f
C208 cp1_buffer1_2/charge_pump1_0/capacitors_1_12/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# cp1_buffer1_2/charge_pump1_0/vdd 13.3f
C209 cp1_buffer1_reverse_0/charge_pump1_reverse_0/capacitor_8_1/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# VSUBS 6.15f
C210 cp1_buffer1_2/charge_pump1_0/in4 cp1_buffer1_2/charge_pump1_0/vdd 13.9f
C211 cp1_buffer1_2/charge_pump1_0/capacitors_1_2/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# cp1_buffer1_2/charge_pump1_0/clk 2.17f
C212 cp1_buffer1_reverse_1/charge_pump1_reverse_0/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# cp1_buffer1_reverse_1/charge_pump1_reverse_0/clock_1/clkb 2.17f
C213 cp1_buffer1_reverse_1/charge_pump1_reverse_0/capacitors_1_10/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# cp1_buffer1_reverse_1/charge_pump1_reverse_0/capacitors_1_10/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/m1_5444_838# 2.1f
C214 cp1_buffer1_0/charge_pump1_0/capacitors_1_13/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# cp1_buffer1_2/charge_pump1_0/vdd 3.48f
C215 cp1_buffer1_2/charge_pump1_0/capacitor_8_1/capacitor_7_0/buffer_and_gate_0/m1_5444_838# cp1_buffer1_2/charge_pump1_0/capacitor_8_1/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 2.1f
C216 cp1_buffer1_2/charge_pump1_0/capacitors_1_11/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# cp1_buffer1_2/charge_pump1_0/vdd 3.49f
C217 VSUBS cp1_buffer1_2/charge_pump1_0/capacitors_1_3/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 6.15f
C218 cp1_buffer1_reverse_0/charge_pump1_reverse_0/capacitors_1_2/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 cp1_buffer1_2/charge_pump1_0/in7 2.94f
C219 cp1_buffer1_2/charge_pump1_0/capacitors_1_5/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/m1_5444_838# cp1_buffer1_2/charge_pump1_0/capacitors_1_5/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 2.1f
C220 VSUBS cp1_buffer1_2/charge_pump1_0/vdd 2p
C221 cp1_buffer1_2/charge_pump1_0/in1 cp1_buffer1_2/charge_pump1_0/capacitors_1_1/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 2.94f
C222 cp1_buffer1_0/charge_pump1_0/clk cp1_buffer1_0/charge_pump1_0/capacitors_1_0/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 2.2f
C223 VSUBS cp1_buffer1_0/charge_pump1_0/input2 10.4f
C224 cp1_buffer1_2/charge_pump1_0/capacitors_1_2/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/m1_5444_838# cp1_buffer1_2/charge_pump1_0/vdd 8.44f
C225 cp1_buffer1_reverse_0/charge_pump1_reverse_0/capacitors_1_13/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/m1_5444_838# VSUBS 4.07f
C226 cp1_buffer1_1/charge_pump1_0/capacitors_1_5/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 cp1_buffer1_2/charge_pump1_0/in3 2.94f
C227 VSUBS cp1_buffer1_1/charge_pump1_0/capacitor_8_1/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 6.15f
C228 cp1_buffer1_2/charge_pump1_0/in3 VSUBS 7.25f
C229 cp1_buffer1_0/charge_pump1_0/clkb cp1_buffer1_0/charge_pump1_0/capacitors_1_1/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 2.18f
C230 cp1_buffer1_0/charge_pump1_0/capacitors_1_0/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/m1_5444_838# cp1_buffer1_2/charge_pump1_0/vdd 8.43f
C231 cp1_buffer1_reverse_0/charge_pump1_reverse_0/clock_1/clk_in cp1_buffer1_2/charge_pump1_0/vdd 9.06f
C232 cp1_buffer1_2/charge_pump1_0/capacitors_1_7/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# cp1_buffer1_2/charge_pump1_0/vdd 3.49f
C233 cp1_buffer1_reverse_1/charge_pump1_reverse_0/capacitors_1_8/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/m1_5444_838# cp1_buffer1_2/charge_pump1_0/vdd 8.44f
C234 cp1_buffer1_2/charge_pump1_0/vdd cp1_buffer1_1/charge_pump1_0/capacitors_1_5/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/m1_5444_838# 8.44f
C235 cp1_buffer1_reverse_1/charge_pump1_reverse_0/capacitors_1_2/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 cp1_buffer1_2/charge_pump1_0/in7 2.94f
C236 cp1_buffer1_reverse_0/charge_pump1_reverse_0/capacitors_1_10/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/m1_5444_838# cp1_buffer1_2/charge_pump1_0/vdd 8.44f
C237 cp1_buffer1_reverse_1/charge_pump1_reverse_0/clock_1/clkb cp1_buffer1_reverse_1/charge_pump1_reverse_0/input1 8.86f
C238 cp1_buffer1_reverse_1/charge_pump1_reverse_0/capacitors_1_8/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# VSUBS 6.15f
C239 cp1_buffer1_1/charge_pump1_0/capacitors_1_12/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# VSUBS 6.15f
C240 cp1_buffer1_reverse_0/charge_pump1_reverse_0/capacitors_1_10/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# VSUBS 6.15f
C241 cp1_buffer1_reverse_1/charge_pump1_reverse_0/capacitors_1_8/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# cp1_buffer1_2/charge_pump1_0/vdd 3.49f
C242 cp1_buffer1_2/charge_pump1_0/vdd cp1_buffer1_0/charge_pump1_0/capacitors_1_9/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 13.3f
C243 cp1_buffer1_reverse_1/charge_pump1_reverse_0/capacitors_1_7/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 cp1_buffer1_2/charge_pump1_0/in4 2.94f
C244 cp1_buffer1_reverse_0/charge_pump1_reverse_0/capacitors_1_10/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# cp1_buffer1_2/charge_pump1_0/vdd 3.48f
C245 cp1_buffer1_2/charge_pump1_0/clk cp1_buffer1_2/charge_pump1_0/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 2.17f
C246 cp1_buffer1_reverse_0/charge_pump1_reverse_0/capacitors_1_8/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/m1_5444_838# VSUBS 4.07f
C247 cp1_buffer1_reverse_0/charge_pump1_reverse_0/clock_1/a_3246_118# cp1_buffer1_2/charge_pump1_0/vdd 7.37f
C248 cp1_buffer1_0/charge_pump1_0/capacitors_1_11/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# cp1_buffer1_2/charge_pump1_0/vdd 13.3f
C249 cp1_buffer1_reverse_1/charge_pump1_reverse_0/capacitors_1_6/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 cp1_buffer1_2/charge_pump1_0/in5 2.94f
C250 cp1_buffer1_2/charge_pump1_0/clk cp1_buffer1_2/charge_pump1_0/capacitors_1_9/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 2.17f
C251 cp1_buffer1_reverse_1/charge_pump1_reverse_0/capacitors_1_12/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# cp1_buffer1_2/charge_pump1_0/vdd 13.3f
C252 VSUBS cp1_buffer1_1/charge_pump1_0/capacitors_1_0/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/m1_5444_838# 4f
C253 cp1_buffer1_reverse_1/charge_pump1_reverse_0/capacitors_1_8/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# cp1_buffer1_reverse_1/charge_pump1_reverse_0/capacitors_1_8/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/m1_5444_838# 2.1f
C254 cp1_buffer1_reverse_1/charge_pump1_reverse_0/clock_1/clkb cp1_buffer1_reverse_1/charge_pump1_reverse_0/clock_1/a_2432_n962# 2.69f
C255 cp1_buffer1_reverse_0/charge_pump1_reverse_0/clock_1/clkb cp1_buffer1_reverse_0/charge_pump1_reverse_0/capacitors_1_9/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 2.17f
C256 cp1_buffer1_1/charge_pump1_0/clk VSUBS 31.6f
C257 cp1_buffer1_reverse_0/charge_pump1_reverse_0/capacitors_1_10/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# cp1_buffer1_reverse_0/charge_pump1_reverse_0/capacitors_1_10/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/m1_5444_838# 2.1f
C258 cp1_buffer1_1/charge_pump1_0/capacitors_1_8/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 cp1_buffer1_2/charge_pump1_0/in6 2.94f
C259 cp1_buffer1_1/charge_pump1_0/capacitors_1_3/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# cp1_buffer1_1/charge_pump1_0/capacitors_1_3/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/m1_5444_838# 2.1f
C260 cp1_buffer1_2/charge_pump1_0/vdd cp1_buffer1_1/charge_pump1_0/capacitors_1_6/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# 3.49f
C261 cp1_buffer1_2/charge_pump1_0/vdd cp1_buffer1_reverse_0/charge_pump1_reverse_0/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/m1_5444_838# 8.43f
C262 cp1_buffer1_0/charge_pump1_0/clkb cp1_buffer1_0/charge_pump1_0/clock_0/a_2432_n962# 2.67f
C263 cp1_buffer1_0/charge_pump1_0/capacitors_1_0/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# cp1_buffer1_2/charge_pump1_0/vdd 13.1f
C264 cp1_buffer1_reverse_0/charge_pump1_reverse_0/input1 VSUBS 9.98f
C265 cp1_buffer1_reverse_0/charge_pump1_reverse_0/capacitors_1_3/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# cp1_buffer1_2/charge_pump1_0/vdd 13.3f
C266 cp1_buffer1_reverse_0/charge_pump1_reverse_0/capacitors_1_7/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# cp1_buffer1_reverse_0/charge_pump1_reverse_0/clock_1/clkb 2.17f
C267 cp1_buffer1_2/charge_pump1_0/vdd cp1_buffer1_2/charge_pump1_0/clock_0/a_2432_n962# 7.04f
C268 cp1_buffer1_reverse_1/charge_pump1_reverse_0/clock_1/clk cp1_buffer1_reverse_1/charge_pump1_reverse_0/capacitors_1_13/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 2.17f
C269 cp1_buffer1_0/charge_pump1_0/capacitors_1_10/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 cp1_buffer1_2/charge_pump1_0/in7 2.94f
C270 cp1_buffer1_reverse_1/charge_pump1_reverse_0/capacitors_1_7/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/m1_5444_838# VSUBS 4.07f
C271 cp1_buffer1_0/charge_pump1_0/capacitors_1_12/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# cp1_buffer1_0/charge_pump1_0/clkb 2.17f
C272 cp1_buffer1_reverse_1/charge_pump1_reverse_0/capacitors_1_2/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# cp1_buffer1_2/charge_pump1_0/vdd 3.49f
C273 cp1_buffer1_2/charge_pump1_0/in4 cp1_buffer1_0/charge_pump1_0/capacitors_1_6/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 2.94f
C274 cp1_buffer1_1/charge_pump1_0/clk cp1_buffer1_1/charge_pump1_0/m1_4341_n519# 9.42f
C275 cp1_buffer1_0/charge_pump1_0/clk cp1_buffer1_0/charge_pump1_0/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 2.17f
C276 cp1_buffer1_0/charge_pump1_0/capacitor_8_1/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# cp1_buffer1_2/charge_pump1_0/vdd 3.48f
C277 VSUBS cp1_buffer1_1/charge_pump1_0/capacitor_8_1/capacitor_7_0/buffer_and_gate_0/m1_5444_838# 4.07f
C278 cp1_buffer1_reverse_1/charge_pump1_reverse_0/capacitors_1_13/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/m1_5444_838# cp1_buffer1_2/charge_pump1_0/vdd 8.43f
C279 cp1_buffer1_2/charge_pump1_0/capacitors_1_8/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# cp1_buffer1_2/charge_pump1_0/capacitors_1_8/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/m1_5444_838# 2.1f
C280 cp1_buffer1_0/charge_pump1_0/capacitors_1_1/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# cp1_buffer1_2/charge_pump1_0/vdd 13.1f
C281 cp1_buffer1_reverse_0/charge_pump1_reverse_0/capacitors_1_4/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/m1_5444_838# VSUBS 4.07f
C282 cp1_buffer1_reverse_0/charge_pump1_reverse_0/capacitors_1_2/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/m1_5444_838# VSUBS 4.07f
C283 cp1_buffer1_2/charge_pump1_0/capacitors_1_8/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 cp1_buffer1_2/charge_pump1_0/in6 2.94f
C284 cp1_buffer1_0/charge_pump1_0/capacitors_1_2/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# VSUBS 6.15f
C285 cp1_buffer1_1/charge_pump1_0/clkb cp1_buffer1_1/charge_pump1_0/capacitors_1_13/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 2.17f
C286 cp1_buffer1_reverse_1/charge_pump1_reverse_0/clock_1/a_2402_572# cp1_buffer1_2/charge_pump1_0/vdd 2.67f
C287 cp1_buffer1_reverse_1/charge_pump1_reverse_0/capacitors_1_13/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# VSUBS 6.15f
C288 cp1_buffer1_0/charge_pump1_0/capacitors_1_10/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# VSUBS 6.15f
C289 cp1_buffer1_0/charge_pump1_0/clk cp1_buffer1_0/charge_pump1_0/capacitors_1_8/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 2.17f
C290 cp1_buffer1_2/charge_pump1_0/capacitors_1_13/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# cp1_buffer1_2/charge_pump1_0/vdd 3.48f
C291 VSUBS cp1_buffer1_2/charge_pump1_0/capacitors_1_1/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 6.05f
C292 VSUBS cp1_buffer1_0/charge_pump1_0/capacitors_1_8/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/m1_5444_838# 4.07f
C293 cp1_buffer1_1/charge_pump1_0/clkb cp1_buffer1_1/charge_pump1_0/capacitors_1_1/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 2.18f
C294 cp1_buffer1_2/charge_pump1_0/capacitors_1_6/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/m1_5444_838# cp1_buffer1_2/charge_pump1_0/vdd 8.43f
C295 cp1_buffer1_reverse_1/charge_pump1_reverse_0/capacitors_1_2/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# cp1_buffer1_2/charge_pump1_0/vdd 13.3f
C296 cp1_buffer1_reverse_1/charge_pump1_reverse_0/capacitors_1_13/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# cp1_buffer1_2/charge_pump1_0/vdd 3.48f
C297 cp1_buffer1_reverse_1/charge_pump1_reverse_0/capacitors_1_6/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# cp1_buffer1_reverse_1/charge_pump1_reverse_0/clock_1/clkb 2.17f
C298 cp1_buffer1_2/charge_pump1_0/in1 cp1_buffer1_1/charge_pump1_0/capacitors_1_1/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 2.94f
C299 cp1_buffer1_2/charge_pump1_0/vdd cp1_buffer1_1/charge_pump1_0/capacitors_1_6/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 13.3f
C300 cp1_buffer1_reverse_1/charge_pump1_reverse_0/clock_1/clkb cp1_buffer1_reverse_1/charge_pump1_reverse_0/capacitors_1_0/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 2.2f
C301 cp1_buffer1_reverse_0/charge_pump1_reverse_0/m1_12659_300# cp1_buffer1_reverse_0/charge_pump1_reverse_0/clock_1/clk 9.24f
C302 cp1_buffer1_2/charge_pump1_0/in5 cp1_buffer1_2/charge_pump1_0/capacitors_1_7/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 2.94f
C303 cp1_buffer1_2/charge_pump1_0/capacitors_1_11/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/m1_5444_838# cp1_buffer1_2/charge_pump1_0/vdd 8.44f
C304 cp1_buffer1_reverse_1/charge_pump1_reverse_0/capacitors_1_1/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/m1_5444_838# VSUBS 4f
C305 cp1_buffer1_2/charge_pump1_0/capacitor_8_1/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# VSUBS 6.15f
C306 cp1_buffer1_1/charge_pump1_0/clkb cp1_buffer1_reverse_1/charge_pump1_reverse_0/nmos_dnw3_0/vs 2.21f
C307 cp1_buffer1_2/charge_pump1_0/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/m1_5444_838# cp1_buffer1_2/charge_pump1_0/vdd 8.43f
C308 cp1_buffer1_reverse_0/charge_pump1_reverse_0/capacitors_1_1/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/m1_5444_838# cp1_buffer1_2/charge_pump1_0/vdd 8.43f
C309 cp1_buffer1_2/charge_pump1_0/clk cp1_buffer1_2/charge_pump1_0/capacitors_1_7/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 2.17f
C310 cp1_buffer1_reverse_1/charge_pump1_reverse_0/capacitors_1_10/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# cp1_buffer1_2/charge_pump1_0/vdd 13.3f
C311 cp1_buffer1_reverse_1/charge_pump1_reverse_0/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# cp1_buffer1_2/charge_pump1_0/vdd 13.3f
C312 cp1_buffer1_2/charge_pump1_0/capacitors_1_0/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/m1_5444_838# cp1_buffer1_2/charge_pump1_0/vdd 8.43f
C313 cp1_buffer1_0/charge_pump1_0/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/m1_5444_838# cp1_buffer1_0/charge_pump1_0/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 2.1f
C314 cp1_buffer1_0/charge_pump1_0/clk cp1_buffer1_0/charge_pump1_0/capacitors_1_3/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 2.17f
C315 cp1_buffer1_reverse_1/charge_pump1_reverse_0/capacitors_1_9/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# cp1_buffer1_2/charge_pump1_0/vdd 3.48f
C316 cp1_buffer1_reverse_0/charge_pump1_reverse_0/capacitors_1_1/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# VSUBS 6.05f
C317 cp1_buffer1_2/charge_pump1_0/vdd cp1_buffer1_1/charge_pump1_0/capacitors_1_8/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 13.3f
C318 cp1_buffer1_reverse_0/charge_pump1_reverse_0/capacitor_8_1/capacitor_7_0/buffer_and_gate_0/m1_5444_838# VSUBS 4.07f
C319 cp1_buffer1_2/charge_pump1_0/in1 VSUBS 6.8f
C320 cp1_buffer1_reverse_1/charge_pump1_reverse_0/capacitors_1_9/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/m1_5444_838# cp1_buffer1_2/charge_pump1_0/vdd 8.44f
C321 cp1_buffer1_1/charge_pump1_0/capacitors_1_4/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/m1_5444_838# cp1_buffer1_2/charge_pump1_0/vdd 8.44f
C322 cp1_buffer1_reverse_0/charge_pump1_reverse_0/capacitors_1_6/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/m1_5444_838# cp1_buffer1_2/charge_pump1_0/vdd 8.44f
C323 cp1_buffer1_reverse_0/charge_pump1_reverse_0/capacitors_1_1/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# cp1_buffer1_2/charge_pump1_0/vdd 3.45f
C324 VSUBS cp1_buffer1_0/charge_pump1_0/capacitors_1_1/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/m1_5444_838# 4f
C325 cp1_buffer1_reverse_1/charge_pump1_reverse_0/capacitors_1_9/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# VSUBS 6.15f
C326 cp1_buffer1_2/charge_pump1_0/in5 cp1_buffer1_0/charge_pump1_0/capacitors_1_7/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 2.94f
C327 cp1_buffer1_reverse_0/charge_pump1_reverse_0/capacitors_1_6/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# VSUBS 6.15f
C328 cp1_buffer1_1/charge_pump1_0/clkb cp1_buffer1_2/charge_pump1_0/vdd 75.1f
C329 cp1_buffer1_2/charge_pump1_0/in4 cp1_buffer1_reverse_0/charge_pump1_reverse_0/capacitors_1_12/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 2.94f
C330 cp1_buffer1_1/charge_pump1_0/capacitors_1_4/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# cp1_buffer1_2/charge_pump1_0/vdd 3.48f
C331 cp1_buffer1_0/charge_pump1_0/capacitors_1_6/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/m1_5444_838# cp1_buffer1_2/charge_pump1_0/vdd 8.43f
C332 cp1_buffer1_reverse_0/charge_pump1_reverse_0/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# VSUBS 6.15f
C333 cp1_buffer1_0/charge_pump1_0/clock_0/a_2432_n962# cp1_buffer1_2/charge_pump1_0/vdd 7.04f
C334 cp1_buffer1_reverse_1/charge_pump1_reverse_0/capacitors_1_11/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/m1_5444_838# VSUBS 4.08f
C335 cp1_buffer1_reverse_0/charge_pump1_reverse_0/capacitors_1_6/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# cp1_buffer1_2/charge_pump1_0/vdd 3.49f
C336 cp1_buffer1_reverse_1/charge_pump1_reverse_0/clock_1/clkb cp1_buffer1_reverse_1/charge_pump1_reverse_0/m1_4341_n519# 9.35f
C337 VSUBS cp1_buffer1_1/charge_pump1_0/capacitors_1_5/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 6.15f
C338 cp1_buffer1_2/charge_pump1_0/in8 cp1_buffer1_reverse_0/charge_pump1_reverse_0/capacitors_1_1/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 2.94f
C339 cp1_buffer1_2/charge_pump1_0/in5 cp1_buffer1_reverse_0/charge_pump1_reverse_0/capacitors_1_13/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 2.94f
C340 cp1_buffer1_0/charge_pump1_0/clkb cp1_buffer1_reverse_0/charge_pump1_reverse_0/nmos_dnw3_0/vs 2.21f
C341 cp1_buffer1_2/charge_pump1_0/capacitors_1_5/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# cp1_buffer1_2/charge_pump1_0/vdd 13.3f
C342 cp1_buffer1_2/charge_pump1_0/clock_0/a_2020_n482# cp1_buffer1_2/charge_pump1_0/vdd 2.66f
C343 cp1_buffer1_1/charge_pump1_0/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# cp1_buffer1_2/charge_pump1_0/vdd 13.3f
C344 cp1_buffer1_2/charge_pump1_0/in8 cp1_buffer1_2/charge_pump1_0/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 2.94f
C345 cp1_buffer1_1/charge_pump1_0/clkb cp1_buffer1_1/charge_pump1_0/capacitor_8_1/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 2.16f
C346 cp1_buffer1_2/charge_pump1_0/vdd cp1_buffer1_0/charge_pump1_0/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 13.3f
C347 cp1_buffer1_1/charge_pump1_0/capacitor_8_1/capacitor_7_0/buffer_and_gate_0/in1 cp1_buffer1_2/charge_pump1_0/in8 2.94f
C348 cp1_buffer1_reverse_1/charge_pump1_reverse_0/input1 cp1_buffer1_2/charge_pump1_0/vdd 27.9f
C349 cp1_buffer1_0/charge_pump1_0/capacitors_1_12/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# cp1_buffer1_2/charge_pump1_0/vdd 13.3f
C350 cp1_buffer1_2/charge_pump1_0/in8 VSUBS 6.61f
C351 cp1_buffer1_2/charge_pump1_0/vdd cp1_buffer1_2/charge_pump1_0/in6 14f
C352 cp1_buffer1_2/charge_pump1_0/vdd cp1_buffer1_1/charge_pump1_0/capacitors_1_10/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# 3.48f
C353 cp1_buffer1_0/charge_pump1_0/clk cp1_buffer1_reverse_0/charge_pump1_reverse_0/nmos_dnw3_0/vs 2.31f
C354 cp1_buffer1_reverse_0/charge_pump1_reverse_0/clock_1/clkb VSUBS 28.4f
C355 cp1_buffer1_1/charge_pump1_0/capacitors_1_0/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# VSUBS 6.05f
C356 cp1_buffer1_0/charge_pump1_0/capacitors_1_8/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# cp1_buffer1_2/charge_pump1_0/vdd 13.3f
C357 cp1_buffer1_reverse_0/charge_pump1_reverse_0/capacitors_1_13/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# cp1_buffer1_reverse_0/charge_pump1_reverse_0/clock_1/clk 2.17f
C358 cp1_buffer1_reverse_1/charge_pump1_reverse_0/capacitors_1_4/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# cp1_buffer1_reverse_1/charge_pump1_reverse_0/clock_1/clk 2.16f
C359 cp1_buffer1_1/charge_pump1_0/clk cp1_buffer1_1/charge_pump1_0/capacitors_1_6/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 2.17f
C360 cp1_buffer1_reverse_0/charge_pump1_reverse_0/nmos_dnw3_0/clkb cp1_buffer1_reverse_0/charge_pump1_reverse_0/clock_1/clk 8.35f
C361 cp1_buffer1_1/charge_pump1_0/capacitors_1_5/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# cp1_buffer1_1/charge_pump1_0/capacitors_1_5/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/m1_5444_838# 2.1f
C362 cp1_buffer1_reverse_0/charge_pump1_reverse_0/capacitors_1_0/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/m1_5444_838# cp1_buffer1_2/charge_pump1_0/vdd 8.43f
C363 cp1_buffer1_1/charge_pump1_0/clkb cp1_buffer1_1/charge_pump1_0/capacitors_1_12/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 2.17f
C364 cp1_buffer1_reverse_1/charge_pump1_reverse_0/capacitor_8_1/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# cp1_buffer1_reverse_1/charge_pump1_reverse_0/clock_1/clk 2.16f
C365 cp1_buffer1_2/charge_pump1_0/input1 cp1_buffer1_2/charge_pump1_0/vdd 28.3f
C366 VSUBS cp1_buffer1_1/charge_pump1_0/capacitors_1_11/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 6.15f
C367 cp1_buffer1_reverse_0/charge_pump1_reverse_0/capacitors_1_8/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# cp1_buffer1_2/charge_pump1_0/vdd 13.3f
C368 cp1_buffer1_2/charge_pump1_0/capacitors_1_9/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/m1_5444_838# cp1_buffer1_2/charge_pump1_0/capacitors_1_9/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 2.1f
C369 cp1_buffer1_2/charge_pump1_0/in8 cp1_buffer1_2/charge_pump1_0/capacitor_8_1/capacitor_7_0/buffer_and_gate_0/in1 2.94f
C370 cp1_buffer1_0/charge_pump1_0/capacitors_1_5/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# cp1_buffer1_0/charge_pump1_0/capacitors_1_5/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/m1_5444_838# 2.1f
C371 cp1_buffer1_reverse_1/charge_pump1_reverse_0/clock_1/clk cp1_buffer1_reverse_1/charge_pump1_reverse_0/clock_1/a_3246_118# 2.73f
C372 cp1_buffer1_reverse_0/charge_pump1_reverse_0/capacitors_1_5/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/m1_5444_838# VSUBS 4.07f
C373 cp1_buffer1_2/charge_pump1_0/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# cp1_buffer1_2/charge_pump1_0/vdd 3.48f
C374 cp1_buffer1_reverse_1/charge_pump1_reverse_0/clock_1/a_2432_n962# cp1_buffer1_2/charge_pump1_0/vdd 7.04f
C375 cp1_buffer1_reverse_0/charge_pump1_reverse_0/capacitors_1_11/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 cp1_buffer1_2/charge_pump1_0/in3 2.94f
C376 cp1_buffer1_reverse_1/charge_pump1_reverse_0/capacitors_1_4/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/m1_5444_838# cp1_buffer1_2/charge_pump1_0/vdd 8.43f
C377 cp1_buffer1_reverse_1/charge_pump1_reverse_0/capacitors_1_0/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 cp1_buffer1_2/charge_pump1_0/in8 2.94f
C378 cp1_buffer1_1/charge_pump1_0/clk cp1_buffer1_1/charge_pump1_0/capacitors_1_8/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 2.17f
C379 cp1_buffer1_reverse_0/charge_pump1_reverse_0/clock_1/a_2402_572# cp1_buffer1_2/charge_pump1_0/vdd 2.67f
C380 cp1_buffer1_2/charge_pump1_0/in5 cp1_buffer1_2/charge_pump1_0/vdd 13.9f
C381 cp1_buffer1_0/charge_pump1_0/clk cp1_buffer1_0/charge_pump1_0/clock_0/a_3246_118# 2.71f
C382 cp1_buffer1_2/charge_pump1_0/vdd cp1_buffer1_0/charge_pump1_0/capacitors_1_3/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 13.3f
C383 cp1_buffer1_1/charge_pump1_0/capacitors_1_10/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 cp1_buffer1_2/charge_pump1_0/in7 2.94f
C384 VSUBS cp1_buffer1_0/charge_pump1_0/capacitors_1_7/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 6.15f
C385 cp1_buffer1_reverse_1/charge_pump1_reverse_0/capacitors_1_13/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# cp1_buffer1_reverse_1/charge_pump1_reverse_0/capacitors_1_13/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/m1_5444_838# 2.1f
C386 cp1_buffer1_2/charge_pump1_0/capacitors_1_10/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# cp1_buffer1_2/charge_pump1_0/clkb 2.16f
C387 cp1_buffer1_reverse_0/charge_pump1_reverse_0/input2 VSUBS 9.75f
C388 cp1_buffer1_reverse_1/charge_pump1_reverse_0/capacitors_1_4/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# VSUBS 6.15f
C389 cp1_buffer1_reverse_1/charge_pump1_reverse_0/capacitors_1_7/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# cp1_buffer1_reverse_1/charge_pump1_reverse_0/clock_1/clkb 2.17f
C390 cp1_buffer1_0/charge_pump1_0/input1 cp1_buffer1_0/charge_pump1_0/clk 8.87f
C391 cp1_buffer1_1/charge_pump1_0/capacitors_1_8/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/m1_5444_838# VSUBS 4.07f
C392 cp1_buffer1_reverse_1/charge_pump1_reverse_0/capacitors_1_4/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# cp1_buffer1_2/charge_pump1_0/vdd 3.48f
C393 cp1_buffer1_reverse_1/charge_pump1_reverse_0/capacitor_8_1/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# VSUBS 6.15f
C394 cp1_buffer1_reverse_1/charge_pump1_reverse_0/capacitor_8_1/capacitor_7_0/buffer_and_gate_0/m1_5444_838# cp1_buffer1_2/charge_pump1_0/vdd 8.43f
C395 cp1_buffer1_2/charge_pump1_0/capacitor_8_1/capacitor_7_0/buffer_and_gate_0/m1_5444_838# VSUBS 4.07f
C396 cp1_buffer1_2/charge_pump1_0/clk cp1_buffer1_2/charge_pump1_0/clock_0/a_3246_118# 2.71f
C397 cp1_buffer1_2/charge_pump1_0/in3 cp1_buffer1_0/charge_pump1_0/capacitors_1_5/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 2.94f
C398 cp1_buffer1_2/charge_pump1_0/capacitors_1_5/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 cp1_buffer1_2/charge_pump1_0/in3 2.94f
C399 VSUBS cp1_buffer1_1/charge_pump1_0/capacitors_1_7/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/m1_5444_838# 4.07f
C400 cp1_buffer1_2/charge_pump1_0/clkb cp1_buffer1_2/charge_pump1_0/m1_12464_n576# 2.21f
C401 cp1_buffer1_reverse_0/charge_pump1_reverse_0/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# cp1_buffer1_reverse_0/charge_pump1_reverse_0/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/m1_5444_838# 2.1f
C402 cp1_buffer1_1/charge_pump1_0/capacitors_1_10/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# VSUBS 6.15f
C403 cp1_buffer1_2/charge_pump1_0/capacitors_1_13/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/m1_5444_838# cp1_buffer1_2/charge_pump1_0/vdd 8.43f
C404 cp1_buffer1_0/charge_pump1_0/capacitors_1_11/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/m1_5444_838# VSUBS 4.08f
C405 cp1_buffer1_1/charge_pump1_0/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# cp1_buffer1_1/charge_pump1_0/clk 2.17f
C406 cp1_buffer1_reverse_0/charge_pump1_reverse_0/capacitors_1_9/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/m1_5444_838# cp1_buffer1_2/charge_pump1_0/vdd 8.44f
C407 VSUBS cp1_buffer1_1/charge_pump1_0/capacitors_1_4/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 6.15f
C408 VSUBS cp1_buffer1_2/charge_pump1_0/capacitors_1_3/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/m1_5444_838# 4.07f
C409 VSUBS cp1_buffer1_2/charge_pump1_0/capacitors_1_13/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 6.15f
C410 cp1_buffer1_reverse_1/charge_pump1_reverse_0/m1_12659_300# cp1_buffer1_2/charge_pump1_0/vin 2.14f
C411 cp1_buffer1_reverse_1/charge_pump1_reverse_0/capacitors_1_6/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# cp1_buffer1_reverse_1/charge_pump1_reverse_0/capacitors_1_6/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/m1_5444_838# 2.1f
C412 cp1_buffer1_2/charge_pump1_0/input2 cp1_buffer1_2/charge_pump1_0/vdd 28f
C413 cp1_buffer1_reverse_0/charge_pump1_reverse_0/capacitors_1_9/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# VSUBS 6.15f
C414 cp1_buffer1_2/charge_pump1_0/capacitors_1_10/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# cp1_buffer1_2/charge_pump1_0/vdd 3.48f
C415 cp1_buffer1_reverse_0/charge_pump1_reverse_0/capacitors_1_7/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/m1_5444_838# cp1_buffer1_2/charge_pump1_0/vdd 8.44f
C416 cp1_buffer1_2/charge_pump1_0/vdd cp1_buffer1_1/charge_pump1_0/capacitors_1_3/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/m1_5444_838# 8.44f
C417 cp1_buffer1_reverse_0/charge_pump1_reverse_0/capacitors_1_8/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# cp1_buffer1_reverse_0/charge_pump1_reverse_0/capacitors_1_8/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/m1_5444_838# 2.1f
C418 cp1_buffer1_reverse_0/charge_pump1_reverse_0/capacitors_1_9/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# cp1_buffer1_2/charge_pump1_0/vdd 3.48f
C419 cp1_buffer1_2/charge_pump1_0/vdd cp1_buffer1_reverse_0/charge_pump1_reverse_0/nmos_dnw3_0/vs 10.6f
C420 cp1_buffer1_1/charge_pump1_0/input1 cp1_buffer1_1/charge_pump1_0/input2 3.33f
C421 cp1_buffer1_reverse_1/charge_pump1_reverse_0/capacitors_1_0/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# cp1_buffer1_2/charge_pump1_0/vdd 3.45f
C422 cp1_buffer1_0/charge_pump1_0/capacitors_1_1/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/m1_5444_838# cp1_buffer1_0/charge_pump1_0/capacitors_1_1/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 2.1f
C423 cp1_buffer1_reverse_0/charge_pump1_reverse_0/capacitors_1_7/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# VSUBS 6.15f
C424 cp1_buffer1_2/charge_pump1_0/capacitors_1_8/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# cp1_buffer1_2/charge_pump1_0/vdd 13.3f
C425 cp1_buffer1_2/charge_pump1_0/capacitors_1_6/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# cp1_buffer1_2/charge_pump1_0/vdd 13.3f
C426 cp1_buffer1_0/charge_pump1_0/capacitors_1_4/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/m1_5444_838# VSUBS 4.07f
C427 VSUBS cp1_buffer1_1/charge_pump1_0/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/m1_5444_838# 4.07f
C428 cp1_buffer1_2/charge_pump1_0/capacitors_1_0/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# VSUBS 6.05f
C429 cp1_buffer1_reverse_1/charge_pump1_reverse_0/capacitors_1_6/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# cp1_buffer1_2/charge_pump1_0/vdd 13.3f
C430 cp1_buffer1_reverse_0/charge_pump1_reverse_0/capacitors_1_3/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# cp1_buffer1_reverse_0/charge_pump1_reverse_0/clock_1/clkb 2.17f
C431 cp1_buffer1_1/charge_pump1_0/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# cp1_buffer1_2/charge_pump1_0/vdd 3.48f
C432 cp1_buffer1_1/charge_pump1_0/capacitors_1_0/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# cp1_buffer1_2/charge_pump1_0/vdd 3.45f
C433 cp1_buffer1_reverse_0/charge_pump1_reverse_0/capacitors_1_7/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# cp1_buffer1_2/charge_pump1_0/vdd 3.49f
C434 cp1_buffer1_2/charge_pump1_0/clk cp1_buffer1_2/charge_pump1_0/m1_12464_n576# 2.31f
C435 cp1_buffer1_2/charge_pump1_0/in2 cp1_buffer1_2/charge_pump1_0/capacitors_1_4/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 2.94f
C436 cp1_buffer1_reverse_1/charge_pump1_reverse_0/capacitors_1_0/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# cp1_buffer1_2/charge_pump1_0/vdd 13.1f
C437 cp1_buffer1_2/charge_pump1_0/capacitors_1_11/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# VSUBS 6.15f
C438 cp1_buffer1_reverse_1/charge_pump1_reverse_0/capacitors_1_3/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/m1_5444_838# VSUBS 4.07f
C439 cp1_buffer1_1/charge_pump1_0/m1_12659_300# cp1_buffer1_reverse_1/charge_pump1_reverse_0/nmos_dnw3_0/vs 2.14f
C440 cp1_buffer1_2/charge_pump1_0/capacitors_1_4/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# VSUBS 6.15f
C441 cp1_buffer1_0/charge_pump1_0/m1_12659_300# cp1_buffer1_reverse_0/charge_pump1_reverse_0/nmos_dnw3_0/vs 2.14f
C442 cp1_buffer1_1/charge_pump1_0/vin cp1_buffer1_2/charge_pump1_0/vdd 10.3f
C443 cp1_buffer1_reverse_0/charge_pump1_reverse_0/capacitors_1_1/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# cp1_buffer1_reverse_0/charge_pump1_reverse_0/capacitors_1_1/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/m1_5444_838# 2.1f
C444 cp1_buffer1_0/charge_pump1_0/capacitors_1_9/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/m1_5444_838# cp1_buffer1_2/charge_pump1_0/vdd 8.44f
C445 cp1_buffer1_1/charge_pump1_0/input2 cp1_buffer1_2/charge_pump1_0/vdd 28f
C446 cp1_buffer1_2/charge_pump1_0/clkb cp1_buffer1_2/charge_pump1_0/vdd 75.2f
C447 cp1_buffer1_0/charge_pump1_0/clock_0/a_3246_118# cp1_buffer1_2/charge_pump1_0/vdd 7.35f
C448 cp1_buffer1_reverse_0/charge_pump1_reverse_0/capacitors_1_13/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# cp1_buffer1_2/charge_pump1_0/vdd 13.3f
C449 cp1_buffer1_2/charge_pump1_0/capacitors_1_6/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# cp1_buffer1_2/charge_pump1_0/vdd 3.49f
C450 cp1_buffer1_reverse_0/charge_pump1_reverse_0/capacitors_1_4/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# cp1_buffer1_reverse_0/charge_pump1_reverse_0/clock_1/clk 2.16f
C451 cp1_buffer1_0/charge_pump1_0/capacitors_1_11/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# cp1_buffer1_0/charge_pump1_0/capacitors_1_11/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/m1_5444_838# 2.1f
C452 cp1_buffer1_0/charge_pump1_0/capacitors_1_3/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/m1_5444_838# cp1_buffer1_2/charge_pump1_0/vdd 8.44f
C453 cp1_buffer1_2/charge_pump1_0/capacitors_1_9/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# cp1_buffer1_2/charge_pump1_0/vdd 3.48f
C454 cp1_buffer1_reverse_1/charge_pump1_reverse_0/capacitors_1_5/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# cp1_buffer1_reverse_1/charge_pump1_reverse_0/clock_1/clk 2.16f
C455 cp1_buffer1_reverse_0/charge_pump1_reverse_0/capacitors_1_13/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# cp1_buffer1_reverse_0/charge_pump1_reverse_0/capacitors_1_13/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/m1_5444_838# 2.1f
C456 cp1_buffer1_reverse_0/charge_pump1_reverse_0/capacitors_1_9/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 cp1_buffer1_2/charge_pump1_0/in2 2.94f
C457 cp1_buffer1_0/charge_pump1_0/input1 cp1_buffer1_2/charge_pump1_0/vdd 28.3f
C458 cp1_buffer1_2/charge_pump1_0/in2 cp1_buffer1_0/charge_pump1_0/capacitors_1_4/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 2.94f
C459 cp1_buffer1_reverse_0/charge_pump1_reverse_0/capacitors_1_4/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 cp1_buffer1_2/charge_pump1_0/in7 2.94f
C460 cp1_buffer1_reverse_1/charge_pump1_reverse_0/capacitors_1_9/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# cp1_buffer1_reverse_1/charge_pump1_reverse_0/capacitors_1_9/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/m1_5444_838# 2.1f
C461 cp1_buffer1_0/charge_pump1_0/capacitors_1_5/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/m1_5444_838# cp1_buffer1_2/charge_pump1_0/vdd 8.44f
C462 cp1_buffer1_2/charge_pump1_0/in2 cp1_buffer1_reverse_1/charge_pump1_reverse_0/capacitors_1_10/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 2.94f
C463 cp1_buffer1_0/charge_pump1_0/input1 cp1_buffer1_0/charge_pump1_0/input2 3.33f
C464 cp1_buffer1_reverse_1/charge_pump1_reverse_0/capacitors_1_0/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/m1_5444_838# VSUBS 4f
C465 cp1_buffer1_0/charge_pump1_0/capacitors_1_8/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# cp1_buffer1_0/charge_pump1_0/capacitors_1_8/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/m1_5444_838# 2.1f
C466 cp1_buffer1_2/charge_pump1_0/m1_12659_300# cp1_buffer1_2/charge_pump1_0/clkb 9.47f
C467 cp1_buffer1_0/charge_pump1_0/capacitors_1_10/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/m1_5444_838# cp1_buffer1_2/charge_pump1_0/vdd 8.44f
C468 cp1_buffer1_1/charge_pump1_0/capacitors_1_9/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/m1_5444_838# cp1_buffer1_1/charge_pump1_0/capacitors_1_9/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 2.1f
C469 cp1_buffer1_reverse_0/charge_pump1_reverse_0/capacitors_1_6/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# cp1_buffer1_reverse_0/charge_pump1_reverse_0/capacitors_1_6/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/m1_5444_838# 2.1f
C470 cp1_buffer1_2/charge_pump1_0/capacitors_1_2/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# cp1_buffer1_2/charge_pump1_0/vdd 13.3f
C471 cp1_buffer1_reverse_1/charge_pump1_reverse_0/capacitors_1_5/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/m1_5444_838# cp1_buffer1_2/charge_pump1_0/vdd 8.44f
C472 cp1_buffer1_reverse_0/charge_pump1_reverse_0/capacitors_1_12/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/m1_5444_838# VSUBS 4.07f
C473 cp1_buffer1_2/charge_pump1_0/clk cp1_buffer1_2/charge_pump1_0/capacitors_1_3/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 2.17f
C474 cp1_buffer1_2/charge_pump1_0/vdd cp1_buffer1_0/charge_pump1_0/capacitors_1_9/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# 3.48f
C475 cp1_buffer1_reverse_1/charge_pump1_reverse_0/input2 cp1_buffer1_2/charge_pump1_0/vdd 28f
C476 cp1_buffer1_2/charge_pump1_0/clk cp1_buffer1_2/charge_pump1_0/vdd 82.4f
C477 cp1_buffer1_reverse_1/charge_pump1_reverse_0/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/m1_5444_838# cp1_buffer1_2/charge_pump1_0/vdd 8.43f
C478 cp1_buffer1_0/charge_pump1_0/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# cp1_buffer1_2/charge_pump1_0/vdd 3.48f
C479 cp1_buffer1_2/charge_pump1_0/in2 cp1_buffer1_0/charge_pump1_0/capacitors_1_2/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 2.94f
C480 cp1_buffer1_reverse_1/charge_pump1_reverse_0/capacitors_1_5/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# VSUBS 6.15f
C481 cp1_buffer1_1/charge_pump1_0/clkb cp1_buffer1_1/charge_pump1_0/capacitors_1_5/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 2.16f
C482 cp1_buffer1_reverse_1/charge_pump1_reverse_0/capacitors_1_5/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# cp1_buffer1_2/charge_pump1_0/vdd 3.48f
C483 cp1_buffer1_2/charge_pump1_0/capacitors_1_7/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/m1_5444_838# VSUBS 4.07f
C484 cp1_buffer1_0/charge_pump1_0/clk_in VSUBS 6.28f
C485 cp1_buffer1_2/charge_pump1_0/vdd cp1_buffer1_2/charge_pump1_0/in7 13.6f
C486 cp1_buffer1_reverse_1/charge_pump1_reverse_0/clock_1/clk VSUBS 30.9f
C487 cp1_buffer1_reverse_0/charge_pump1_reverse_0/capacitors_1_11/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/m1_5444_838# cp1_buffer1_2/charge_pump1_0/vdd 8.44f
C488 cp1_buffer1_0/charge_pump1_0/capacitors_1_6/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# cp1_buffer1_2/charge_pump1_0/vdd 3.49f
C489 cp1_buffer1_1/charge_pump1_0/capacitors_1_2/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/m1_5444_838# cp1_buffer1_1/charge_pump1_0/capacitors_1_2/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 2.1f
C490 cp1_buffer1_reverse_0/charge_pump1_reverse_0/capacitors_1_0/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# cp1_buffer1_2/charge_pump1_0/vdd 13.1f
C491 cp1_buffer1_2/charge_pump1_0/capacitors_1_12/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/m1_5444_838# cp1_buffer1_2/charge_pump1_0/vdd 8.44f
C492 cp1_buffer1_0/charge_pump1_0/capacitors_1_6/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# VSUBS 6.15f
C493 cp1_buffer1_2/charge_pump1_0/vdd cp1_buffer1_0/charge_pump1_0/capacitors_1_12/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/m1_5444_838# 8.44f
C494 cp1_buffer1_reverse_0/charge_pump1_reverse_0/capacitors_1_11/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# VSUBS 6.15f
C495 cp1_buffer1_1/charge_pump1_0/capacitors_1_6/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/m1_5444_838# VSUBS 4.07f
C496 cp1_buffer1_1/charge_pump1_0/vin cp1_buffer1_1/charge_pump1_0/clk 2.19f
C497 cp1_buffer1_1/charge_pump1_0/capacitors_1_1/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/m1_5444_838# cp1_buffer1_1/charge_pump1_0/capacitors_1_1/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 2.1f
C498 cp1_buffer1_2/charge_pump1_0/capacitors_1_12/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# VSUBS 6.15f
C499 cp1_buffer1_reverse_0/charge_pump1_reverse_0/capacitors_1_11/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# cp1_buffer1_2/charge_pump1_0/vdd 3.49f
C500 cp1_buffer1_2/charge_pump1_0/in4 VSUBS 7.29f
C501 cp1_buffer1_reverse_0/charge_pump1_reverse_0/capacitors_1_5/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 cp1_buffer1_2/charge_pump1_0/in6 2.94f
C502 cp1_buffer1_2/charge_pump1_0/in8 cp1_buffer1_reverse_1/charge_pump1_reverse_0/capacitors_1_1/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 2.94f
C503 cp1_buffer1_1/charge_pump1_0/clkb cp1_buffer1_1/charge_pump1_0/capacitors_1_11/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 2.16f
C504 cp1_buffer1_2/charge_pump1_0/capacitors_1_3/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# cp1_buffer1_2/charge_pump1_0/vdd 3.48f
C505 cp1_buffer1_2/charge_pump1_0/vin cp1_buffer1_2/charge_pump1_0/clk 2.19f
C506 cp1_buffer1_1/charge_pump1_0/capacitors_1_11/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 cp1_buffer1_2/charge_pump1_0/in6 2.94f
C507 cp1_buffer1_2/charge_pump1_0/capacitors_1_10/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# cp1_buffer1_2/charge_pump1_0/capacitors_1_10/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/m1_5444_838# 2.1f
C508 cp1_buffer1_reverse_1/charge_pump1_reverse_0/capacitors_1_7/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# cp1_buffer1_2/charge_pump1_0/vdd 13.3f
C509 cp1_buffer1_0/charge_pump1_0/clk cp1_buffer1_0/charge_pump1_0/vin 2.19f
C510 cp1_buffer1_1/charge_pump1_0/capacitors_1_8/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/m1_5444_838# cp1_buffer1_1/charge_pump1_0/capacitors_1_8/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 2.1f
C511 cp1_buffer1_0/charge_pump1_0/capacitor_8_1/capacitor_7_0/buffer_and_gate_0/m1_5444_838# cp1_buffer1_0/charge_pump1_0/capacitor_8_1/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 2.1f
C512 cp1_buffer1_2/charge_pump1_0/vdd cp1_buffer1_2/charge_pump1_0/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 13.3f
C513 cp1_buffer1_2/charge_pump1_0/capacitors_1_2/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/m1_5444_838# VSUBS 4.07f
C514 cp1_buffer1_2/charge_pump1_0/capacitors_1_9/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# cp1_buffer1_2/charge_pump1_0/vdd 13.3f
C515 cp1_buffer1_1/charge_pump1_0/capacitors_1_12/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/m1_5444_838# cp1_buffer1_2/charge_pump1_0/vdd 8.44f
C516 cp1_buffer1_0/charge_pump1_0/capacitors_1_0/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/m1_5444_838# VSUBS 4f
C517 cp1_buffer1_reverse_0/charge_pump1_reverse_0/clock_1/clk_in VSUBS 5.97f
C518 cp1_buffer1_reverse_0/charge_pump1_reverse_0/capacitors_1_4/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# cp1_buffer1_2/charge_pump1_0/vdd 13.3f
C519 cp1_buffer1_2/charge_pump1_0/in7 cp1_buffer1_1/charge_pump1_0/capacitors_1_9/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 2.94f
C520 cp1_buffer1_reverse_0/charge_pump1_reverse_0/capacitors_1_8/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# cp1_buffer1_reverse_0/charge_pump1_reverse_0/clock_1/clkb 2.17f
C521 cp1_buffer1_reverse_0/charge_pump1_reverse_0/capacitors_1_2/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# cp1_buffer1_2/charge_pump1_0/vdd 13.3f
C522 cp1_buffer1_1/charge_pump1_0/capacitors_1_4/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/m1_5444_838# cp1_buffer1_1/charge_pump1_0/capacitors_1_4/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 2.1f
C523 cp1_buffer1_reverse_0/charge_pump1_reverse_0/capacitors_1_5/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# cp1_buffer1_reverse_0/charge_pump1_reverse_0/clock_1/clk 2.16f
C524 cp1_buffer1_reverse_1/charge_pump1_reverse_0/clock_1/clk cp1_buffer1_reverse_1/charge_pump1_reverse_0/capacitors_1_12/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 2.17f
C525 cp1_buffer1_reverse_1/charge_pump1_reverse_0/capacitors_1_8/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/m1_5444_838# VSUBS 4.07f
C526 cp1_buffer1_1/charge_pump1_0/capacitors_1_1/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/m1_5444_838# cp1_buffer1_2/charge_pump1_0/vdd 8.43f
C527 cp1_buffer1_2/charge_pump1_0/in2 cp1_buffer1_2/charge_pump1_0/vdd 13.9f
C528 VSUBS cp1_buffer1_1/charge_pump1_0/capacitors_1_5/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/m1_5444_838# 4.07f
C529 cp1_buffer1_1/charge_pump1_0/capacitors_1_10/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# cp1_buffer1_1/charge_pump1_0/clkb 2.16f
C530 cp1_buffer1_reverse_0/charge_pump1_reverse_0/capacitors_1_10/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/m1_5444_838# VSUBS 4.07f
C531 cp1_buffer1_2/charge_pump1_0/in1 cp1_buffer1_0/charge_pump1_0/capacitors_1_1/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 2.94f
C532 cp1_buffer1_0/charge_pump1_0/capacitors_1_11/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# cp1_buffer1_2/charge_pump1_0/vdd 3.49f
C533 cp1_buffer1_1/charge_pump1_0/capacitors_1_11/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/m1_5444_838# cp1_buffer1_2/charge_pump1_0/vdd 8.44f
C534 cp1_buffer1_2/charge_pump1_0/vdd cp1_buffer1_1/charge_pump1_0/capacitors_1_9/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 13.3f
C535 cp1_buffer1_2/charge_pump1_0/capacitors_1_0/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/m1_5444_838# cp1_buffer1_2/charge_pump1_0/capacitors_1_0/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 2.1f
C536 cp1_buffer1_2/charge_pump1_0/clkb cp1_buffer1_2/charge_pump1_0/capacitors_1_1/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 2.18f
C537 cp1_buffer1_1/charge_pump1_0/clkb cp1_buffer1_1/charge_pump1_0/capacitors_1_4/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 2.16f
C538 cp1_buffer1_2/charge_pump1_0/capacitors_1_11/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# cp1_buffer1_2/charge_pump1_0/capacitors_1_11/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/m1_5444_838# 2.1f
C539 cp1_buffer1_reverse_1/charge_pump1_reverse_0/capacitors_1_3/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# cp1_buffer1_reverse_1/charge_pump1_reverse_0/clock_1/clkb 2.17f
C540 cp1_buffer1_0/charge_pump1_0/capacitor_8_1/capacitor_7_0/buffer_and_gate_0/m1_5444_838# cp1_buffer1_2/charge_pump1_0/vdd 8.43f
C541 VSUBS cp1_buffer1_0/charge_pump1_0/capacitors_1_9/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 6.15f
C542 cp1_buffer1_reverse_1/charge_pump1_reverse_0/capacitors_1_12/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/m1_5444_838# cp1_buffer1_2/charge_pump1_0/vdd 8.44f
C543 cp1_buffer1_1/charge_pump1_0/capacitors_1_10/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/m1_5444_838# cp1_buffer1_2/charge_pump1_0/vdd 8.44f
C544 cp1_buffer1_reverse_1/charge_pump1_reverse_0/capacitors_1_1/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# cp1_buffer1_2/charge_pump1_0/vdd 13.1f
C545 cp1_buffer1_1/charge_pump1_0/capacitors_1_12/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/m1_5444_838# cp1_buffer1_1/charge_pump1_0/capacitors_1_12/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 2.1f
C546 cp1_buffer1_0/charge_pump1_0/capacitors_1_10/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/m1_5444_838# cp1_buffer1_0/charge_pump1_0/capacitors_1_10/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 2.1f
C547 cp1_buffer1_0/charge_pump1_0/capacitors_1_11/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# VSUBS 6.15f
C548 cp1_buffer1_2/charge_pump1_0/capacitor_8_1/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# cp1_buffer1_2/charge_pump1_0/clkb 2.16f
C549 cp1_buffer1_reverse_1/charge_pump1_reverse_0/capacitors_1_12/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# VSUBS 6.15f
C550 cp1_buffer1_1/charge_pump1_0/capacitors_1_5/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# cp1_buffer1_2/charge_pump1_0/vdd 3.48f
C551 cp1_buffer1_reverse_1/charge_pump1_reverse_0/capacitor_8_1/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# cp1_buffer1_2/charge_pump1_0/vdd 3.48f
C552 cp1_buffer1_reverse_1/charge_pump1_reverse_0/capacitors_1_12/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# cp1_buffer1_2/charge_pump1_0/vdd 3.48f
C553 cp1_buffer1_1/charge_pump1_0/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# cp1_buffer1_1/charge_pump1_0/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/m1_5444_838# 2.1f
C554 cp1_buffer1_reverse_1/charge_pump1_reverse_0/capacitors_1_4/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# cp1_buffer1_reverse_1/charge_pump1_reverse_0/capacitors_1_4/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/m1_5444_838# 2.1f
C555 cp1_buffer1_reverse_0/charge_pump1_reverse_0/capacitors_1_8/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 cp1_buffer1_2/charge_pump1_0/in3 2.94f
C556 cp1_buffer1_2/charge_pump1_0/capacitors_1_10/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/m1_5444_838# cp1_buffer1_2/charge_pump1_0/vdd 8.44f
C557 cp1_buffer1_reverse_0/charge_pump1_reverse_0/capacitors_1_3/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/m1_5444_838# cp1_buffer1_2/charge_pump1_0/vdd 8.44f
C558 cp1_buffer1_2/charge_pump1_0/vdd cp1_buffer1_1/charge_pump1_0/capacitors_1_7/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 13.3f
C559 VSUBS cp1_buffer1_reverse_0/charge_pump1_reverse_0/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/m1_5444_838# 4.07f
C560 cp1_buffer1_0/charge_pump1_0/vin cp1_buffer1_2/charge_pump1_0/vdd 9.13f
C561 cp1_buffer1_reverse_0/charge_pump1_reverse_0/clock_1/clkb cp1_buffer1_reverse_0/charge_pump1_reverse_0/nmos_dnw3_0/vs 2.22f
C562 VSUBS cp1_buffer1_0/charge_pump1_0/capacitors_1_0/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 6.05f
C563 cp1_buffer1_reverse_0/charge_pump1_reverse_0/clock_1/clkb cp1_buffer1_reverse_0/charge_pump1_reverse_0/nmos_dnw3_0/clk 8.37f
C564 cp1_buffer1_1/charge_pump1_0/clkb cp1_buffer1_1/charge_pump1_0/clock_0/a_2432_n962# 2.67f
C565 cp1_buffer1_reverse_1/charge_pump1_reverse_0/capacitors_1_11/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# cp1_buffer1_2/charge_pump1_0/vdd 13.3f
C566 cp1_buffer1_reverse_0/charge_pump1_reverse_0/capacitors_1_3/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# VSUBS 6.15f
C567 cp1_buffer1_1/charge_pump1_0/capacitors_1_13/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/m1_5444_838# cp1_buffer1_1/charge_pump1_0/capacitors_1_13/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 2.1f
C568 cp1_buffer1_reverse_0/charge_pump1_reverse_0/capacitors_1_3/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# cp1_buffer1_2/charge_pump1_0/vdd 3.48f
C569 cp1_buffer1_reverse_1/charge_pump1_reverse_0/capacitors_1_7/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# cp1_buffer1_reverse_1/charge_pump1_reverse_0/capacitors_1_7/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/m1_5444_838# 2.1f
C570 cp1_buffer1_reverse_1/charge_pump1_reverse_0/capacitor_8_1/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# cp1_buffer1_reverse_1/charge_pump1_reverse_0/capacitor_8_1/capacitor_7_0/buffer_and_gate_0/m1_5444_838# 2.1f
C571 cp1_buffer1_0/charge_pump1_0/capacitors_1_5/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# cp1_buffer1_0/charge_pump1_0/clkb 2.16f
C572 cp1_buffer1_1/charge_pump1_0/capacitors_1_3/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 cp1_buffer1_2/charge_pump1_0/in3 2.94f
C573 cp1_buffer1_2/charge_pump1_0/capacitors_1_7/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# cp1_buffer1_2/charge_pump1_0/vdd 13.3f
C574 cp1_buffer1_2/charge_pump1_0/vdd cp1_buffer1_1/charge_pump1_0/capacitors_1_2/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 13.3f
C575 cp1_buffer1_1/charge_pump1_0/capacitors_1_3/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# cp1_buffer1_2/charge_pump1_0/vdd 13.3f
C576 cp1_buffer1_0/charge_pump1_0/capacitors_1_0/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/m1_5444_838# cp1_buffer1_0/charge_pump1_0/capacitors_1_0/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 2.1f
C577 cp1_buffer1_reverse_0/charge_pump1_reverse_0/clock_1/clkb cp1_buffer1_1/charge_pump1_0/vin 2.02f
C578 cp1_buffer1_2/charge_pump1_0/capacitors_1_9/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/m1_5444_838# cp1_buffer1_2/charge_pump1_0/vdd 8.44f
C579 cp1_buffer1_reverse_1/charge_pump1_reverse_0/clock_1/clkb cp1_buffer1_reverse_1/charge_pump1_reverse_0/nmos_dnw3_0/vs 2.22f
C580 cp1_buffer1_1/charge_pump1_0/clk cp1_buffer1_1/charge_pump1_0/capacitors_1_9/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 2.17f
C581 cp1_buffer1_1/charge_pump1_0/capacitors_1_6/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/m1_5444_838# cp1_buffer1_1/charge_pump1_0/capacitors_1_6/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 2.1f
C582 cp1_buffer1_2/charge_pump1_0/capacitors_1_5/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/m1_5444_838# cp1_buffer1_2/charge_pump1_0/vdd 8.44f
C583 cp1_buffer1_reverse_1/charge_pump1_reverse_0/capacitors_1_13/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/m1_5444_838# VSUBS 4.07f
C584 cp1_buffer1_0/charge_pump1_0/capacitors_1_13/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# cp1_buffer1_0/charge_pump1_0/clkb 2.17f
C585 VSUBS cp1_buffer1_0/charge_pump1_0/capacitors_1_1/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 6.05f
C586 cp1_buffer1_2/charge_pump1_0/in8 cp1_buffer1_1/charge_pump1_0/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 2.94f
C587 cp1_buffer1_reverse_1/charge_pump1_reverse_0/clock_1/clk cp1_buffer1_reverse_1/charge_pump1_reverse_0/capacitors_1_10/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 2.16f
C588 cp1_buffer1_reverse_1/charge_pump1_reverse_0/capacitors_1_2/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/m1_5444_838# cp1_buffer1_2/charge_pump1_0/vdd 8.44f
C589 cp1_buffer1_2/charge_pump1_0/in5 cp1_buffer1_2/charge_pump1_0/capacitors_1_12/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 2.94f
C590 cp1_buffer1_2/charge_pump1_0/in1 cp1_buffer1_reverse_0/charge_pump1_reverse_0/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 2.94f
C591 cp1_buffer1_2/charge_pump1_0/capacitors_1_8/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/m1_5444_838# cp1_buffer1_2/charge_pump1_0/vdd 8.44f
C592 cp1_buffer1_2/charge_pump1_0/capacitors_1_13/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# cp1_buffer1_2/charge_pump1_0/capacitors_1_13/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/m1_5444_838# 2.1f
C593 cp1_buffer1_2/charge_pump1_0/capacitors_1_6/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/m1_5444_838# VSUBS 4.07f
C594 cp1_buffer1_reverse_1/charge_pump1_reverse_0/capacitors_1_2/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# VSUBS 6.15f
C595 cp1_buffer1_2/charge_pump1_0/vdd cp1_buffer1_1/charge_pump1_0/capacitors_1_2/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# 3.49f
C596 cp1_buffer1_reverse_0/charge_pump1_reverse_0/capacitors_1_5/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# cp1_buffer1_2/charge_pump1_0/vdd 13.3f
C597 VSUBS cp1_buffer1_1/charge_pump1_0/capacitors_1_6/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 6.15f
C598 cp1_buffer1_reverse_0/charge_pump1_reverse_0/capacitors_1_9/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# cp1_buffer1_reverse_0/charge_pump1_reverse_0/capacitors_1_9/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/m1_5444_838# 2.1f
C599 cp1_buffer1_reverse_0/charge_pump1_reverse_0/capacitors_1_4/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# cp1_buffer1_reverse_0/charge_pump1_reverse_0/capacitors_1_4/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/m1_5444_838# 2.1f
C600 cp1_buffer1_reverse_1/charge_pump1_reverse_0/clock_1/clkb cp1_buffer1_2/charge_pump1_0/vdd 83.5f
C601 cp1_buffer1_reverse_0/charge_pump1_reverse_0/capacitors_1_2/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# cp1_buffer1_reverse_0/charge_pump1_reverse_0/capacitors_1_2/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/m1_5444_838# 2.1f
C602 cp1_buffer1_reverse_1/charge_pump1_reverse_0/capacitors_1_10/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/m1_5444_838# cp1_buffer1_2/charge_pump1_0/vdd 8.44f
C603 cp1_buffer1_reverse_1/charge_pump1_reverse_0/clock_1/clkb cp1_buffer1_reverse_1/charge_pump1_reverse_0/nmos_dnw3_0/clk 8.37f
C604 cp1_buffer1_1/charge_pump1_0/capacitors_1_13/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/m1_5444_838# cp1_buffer1_2/charge_pump1_0/vdd 8.43f
C605 cp1_buffer1_reverse_0/charge_pump1_reverse_0/capacitors_1_12/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# cp1_buffer1_reverse_0/charge_pump1_reverse_0/clock_1/clk 2.17f
C606 cp1_buffer1_reverse_0/charge_pump1_reverse_0/capacitor_8_1/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# cp1_buffer1_2/charge_pump1_0/vdd 3.48f
C607 cp1_buffer1_reverse_1/charge_pump1_reverse_0/capacitors_1_3/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 cp1_buffer1_2/charge_pump1_0/in6 2.94f
C608 cp1_buffer1_2/charge_pump1_0/capacitors_1_11/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/m1_5444_838# VSUBS 4.08f
C609 cp1_buffer1_0/charge_pump1_0/capacitors_1_2/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/m1_5444_838# cp1_buffer1_2/charge_pump1_0/vdd 8.44f
C610 cp1_buffer1_reverse_0/charge_pump1_reverse_0/capacitors_1_1/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/m1_5444_838# VSUBS 4f
C611 cp1_buffer1_2/charge_pump1_0/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/m1_5444_838# VSUBS 4.07f
C612 cp1_buffer1_reverse_1/charge_pump1_reverse_0/capacitors_1_10/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# VSUBS 6.15f
C613 cp1_buffer1_reverse_1/charge_pump1_reverse_0/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# VSUBS 6.15f
C614 cp1_buffer1_2/charge_pump1_0/capacitors_1_0/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/m1_5444_838# VSUBS 4f
C615 cp1_buffer1_0/charge_pump1_0/capacitors_1_1/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# cp1_buffer1_2/charge_pump1_0/vdd 3.45f
C616 cp1_buffer1_1/charge_pump1_0/clk cp1_buffer1_1/charge_pump1_0/capacitors_1_7/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 2.17f
C617 cp1_buffer1_2/charge_pump1_0/clk_in cp1_buffer1_2/charge_pump1_0/vdd 4.45f
C618 cp1_buffer1_0/charge_pump1_0/capacitors_1_6/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/m1_5444_838# cp1_buffer1_0/charge_pump1_0/capacitors_1_6/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 2.1f
C619 cp1_buffer1_reverse_1/charge_pump1_reverse_0/capacitors_1_10/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# cp1_buffer1_2/charge_pump1_0/vdd 3.48f
C620 VSUBS cp1_buffer1_1/charge_pump1_0/capacitors_1_8/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 6.15f
C621 cp1_buffer1_0/charge_pump1_0/clkb cp1_buffer1_0/charge_pump1_0/capacitor_8_1/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 2.16f
C622 cp1_buffer1_reverse_1/charge_pump1_reverse_0/capacitors_1_9/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/m1_5444_838# VSUBS 4.07f
C623 VSUBS cp1_buffer1_1/charge_pump1_0/capacitors_1_4/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/m1_5444_838# 4.07f
C624 cp1_buffer1_reverse_0/charge_pump1_reverse_0/capacitors_1_7/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# cp1_buffer1_reverse_0/charge_pump1_reverse_0/capacitors_1_7/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/m1_5444_838# 2.1f
C625 cp1_buffer1_1/charge_pump1_0/clk_in cp1_buffer1_2/charge_pump1_0/vdd 7.73f
C626 cp1_buffer1_reverse_0/charge_pump1_reverse_0/capacitors_1_6/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/m1_5444_838# VSUBS 4.07f
C627 cp1_buffer1_2/charge_pump1_0/in5 cp1_buffer1_0/charge_pump1_0/capacitors_1_12/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 2.94f
C628 cp1_buffer1_2/charge_pump1_0/in4 cp1_buffer1_0/charge_pump1_0/capacitors_1_13/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 2.94f
C629 cp1_buffer1_2/charge_pump1_0/in8 cp1_buffer1_0/charge_pump1_0/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 2.94f
C630 cp1_buffer1_0/charge_pump1_0/clkb cp1_buffer1_0/charge_pump1_0/capacitors_1_4/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 2.16f
C631 cp1_buffer1_1/charge_pump1_0/clk cp1_buffer1_1/charge_pump1_0/capacitors_1_2/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 2.17f
C632 cp1_buffer1_2/charge_pump1_0/vdd cp1_buffer1_0/charge_pump1_0/capacitors_1_7/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# 3.49f
C633 cp1_buffer1_1/charge_pump1_0/capacitors_1_3/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# cp1_buffer1_1/charge_pump1_0/clk 2.17f
C634 cp1_buffer1_1/charge_pump1_0/capacitors_1_2/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/m1_5444_838# cp1_buffer1_2/charge_pump1_0/vdd 8.44f
C635 cp1_buffer1_1/charge_pump1_0/clkb VSUBS 27.7f
C636 cp1_buffer1_0/charge_pump1_0/capacitors_1_9/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 cp1_buffer1_2/charge_pump1_0/in7 2.94f
C637 cp1_buffer1_0/charge_pump1_0/capacitors_1_13/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/m1_5444_838# cp1_buffer1_0/charge_pump1_0/capacitors_1_13/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 2.1f
C638 cp1_buffer1_reverse_0/charge_pump1_reverse_0/clock_1/clkb cp1_buffer1_reverse_0/charge_pump1_reverse_0/capacitors_1_0/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 2.2f
C639 cp1_buffer1_reverse_0/charge_pump1_reverse_0/capacitor_8_1/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# cp1_buffer1_reverse_0/charge_pump1_reverse_0/clock_1/clk 2.16f
C640 cp1_buffer1_reverse_1/charge_pump1_reverse_0/capacitors_1_8/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# cp1_buffer1_reverse_1/charge_pump1_reverse_0/clock_1/clkb 2.17f
C641 cp1_buffer1_0/charge_pump1_0/capacitors_1_6/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/m1_5444_838# VSUBS 4.07f
C642 cp1_buffer1_2/charge_pump1_0/clkb cp1_buffer1_2/charge_pump1_0/capacitors_1_13/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 2.17f
C643 cp1_buffer1_2/charge_pump1_0/capacitors_1_5/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# VSUBS 6.15f
C644 cp1_buffer1_1/charge_pump1_0/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# VSUBS 6.15f
C645 VSUBS cp1_buffer1_0/charge_pump1_0/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 6.15f
C646 cp1_buffer1_reverse_1/charge_pump1_reverse_0/m1_12659_300# cp1_buffer1_reverse_1/charge_pump1_reverse_0/clock_1/clk 9.24f
C647 cp1_buffer1_reverse_1/charge_pump1_reverse_0/clock_1/clkb cp1_buffer1_2/charge_pump1_0/vin 2.02f
C648 cp1_buffer1_2/charge_pump1_0/vdd cp1_buffer1_reverse_0/charge_pump1_reverse_0/clock_1/clk 78.7f
C649 cp1_buffer1_reverse_1/charge_pump1_reverse_0/input1 VSUBS 9.98f
C650 cp1_buffer1_0/charge_pump1_0/capacitors_1_12/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# VSUBS 6.15f
C651 cp1_buffer1_0/charge_pump1_0/capacitors_1_5/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# cp1_buffer1_2/charge_pump1_0/vdd 13.3f
C652 VSUBS cp1_buffer1_2/charge_pump1_0/in6 7.43f
C653 cp1_buffer1_2/charge_pump1_0/in8 cp1_buffer1_reverse_0/charge_pump1_reverse_0/capacitors_1_0/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 2.94f
C654 cp1_buffer1_2/charge_pump1_0/vdd cp1_buffer1_1/charge_pump1_0/capacitors_1_9/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/m1_5444_838# 8.44f
C655 cp1_buffer1_2/charge_pump1_0/capacitors_1_4/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/m1_5444_838# cp1_buffer1_2/charge_pump1_0/vdd 8.44f
C656 cp1_buffer1_2/charge_pump1_0/vdd cp1_buffer1_2/charge_pump1_0/clock_0/a_3246_118# 7.35f
C657 cp1_buffer1_reverse_1/charge_pump1_reverse_0/capacitors_1_1/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# cp1_buffer1_reverse_1/charge_pump1_reverse_0/capacitors_1_1/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/m1_5444_838# 2.1f
C658 cp1_buffer1_0/charge_pump1_0/clkb cp1_buffer1_2/charge_pump1_0/vdd 75.1f
C659 cp1_buffer1_reverse_1/charge_pump1_reverse_0/capacitors_1_3/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# cp1_buffer1_2/charge_pump1_0/vdd 13.3f
C660 cp1_buffer1_0/charge_pump1_0/capacitors_1_3/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 cp1_buffer1_2/charge_pump1_0/in3 2.94f
C661 cp1_buffer1_0/charge_pump1_0/clkb cp1_buffer1_0/charge_pump1_0/input2 8.93f
C662 cp1_buffer1_0/charge_pump1_0/capacitors_1_8/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# VSUBS 6.15f
C663 cp1_buffer1_2/charge_pump1_0/capacitors_1_11/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# cp1_buffer1_2/charge_pump1_0/clkb 2.16f
C664 cp1_buffer1_0/charge_pump1_0/g2 cp1_buffer1_0/charge_pump1_0/clkb 8.12f
C665 cp1_buffer1_0/charge_pump1_0/capacitors_1_13/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# cp1_buffer1_2/charge_pump1_0/vdd 13.3f
C666 cp1_buffer1_reverse_0/charge_pump1_reverse_0/capacitors_1_0/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/m1_5444_838# VSUBS 4f
C667 cp1_buffer1_reverse_1/charge_pump1_reverse_0/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 cp1_buffer1_2/charge_pump1_0/in1 2.94f
C668 cp1_buffer1_2/charge_pump1_0/capacitors_1_4/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# cp1_buffer1_2/charge_pump1_0/clkb 2.16f
C669 cp1_buffer1_2/charge_pump1_0/input1 VSUBS 9.98f
C670 cp1_buffer1_0/charge_pump1_0/capacitors_1_3/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# cp1_buffer1_2/charge_pump1_0/vdd 3.48f
C671 cp1_buffer1_0/charge_pump1_0/clk cp1_buffer1_2/charge_pump1_0/vdd 82.5f
C672 cp1_buffer1_reverse_0/charge_pump1_reverse_0/capacitors_1_8/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# VSUBS 6.15f
C673 cp1_buffer1_reverse_1/charge_pump1_reverse_0/capacitors_1_0/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# cp1_buffer1_reverse_1/charge_pump1_reverse_0/capacitors_1_0/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/m1_5444_838# 2.1f
C674 cp1_buffer1_2/charge_pump1_0/capacitors_1_10/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# cp1_buffer1_2/charge_pump1_0/vdd 13.3f
C675 cp1_buffer1_reverse_0/charge_pump1_reverse_0/capacitors_1_2/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# cp1_buffer1_reverse_0/charge_pump1_reverse_0/clock_1/clkb 2.17f
C676 cp1_buffer1_0/charge_pump1_0/clkb cp1_buffer1_0/charge_pump1_0/m1_12659_300# 9.47f
C677 cp1_buffer1_reverse_0/charge_pump1_reverse_0/capacitors_1_8/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# cp1_buffer1_2/charge_pump1_0/vdd 3.49f
C678 cp1_buffer1_0/charge_pump1_0/capacitors_1_11/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 cp1_buffer1_2/charge_pump1_0/in6 2.94f
C679 cp1_buffer1_2/charge_pump1_0/in4 cp1_buffer1_reverse_0/charge_pump1_reverse_0/capacitors_1_7/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 2.94f
C680 cp1_buffer1_reverse_1/charge_pump1_reverse_0/capacitors_1_4/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/m1_5444_838# VSUBS 4.07f
C681 cp1_buffer1_reverse_0/charge_pump1_reverse_0/capacitors_1_10/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# cp1_buffer1_reverse_0/charge_pump1_reverse_0/clock_1/clk 2.16f
C682 cp1_buffer1_2/charge_pump1_0/in5 VSUBS 7.23f
C683 VSUBS cp1_buffer1_0/charge_pump1_0/capacitors_1_3/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 6.15f
C684 cp1_buffer1_1/charge_pump1_0/capacitor_8_1/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# cp1_buffer1_2/charge_pump1_0/vdd 3.48f
C685 cp1_buffer1_2/charge_pump1_0/capacitors_1_0/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# cp1_buffer1_2/charge_pump1_0/clk 2.2f
C686 cp1_buffer1_2/charge_pump1_0/vdd cp1_buffer1_0/charge_pump1_0/capacitors_1_7/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/m1_5444_838# 8.44f
C687 cp1_buffer1_reverse_1/charge_pump1_reverse_0/clock_1/clk_in cp1_buffer1_2/charge_pump1_0/vdd 5.99f
C688 cp1_buffer1_reverse_0/charge_pump1_reverse_0/capacitors_1_6/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 cp1_buffer1_2/charge_pump1_0/in5 2.94f
C689 cp1_buffer1_2/charge_pump1_0/vdd cp1_buffer1_1/charge_pump1_0/capacitors_1_13/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 13.3f
C690 cp1_buffer1_reverse_0/charge_pump1_reverse_0/clock_1/clkb cp1_buffer1_reverse_0/charge_pump1_reverse_0/m1_4341_n519# 9.35f
C691 cp1_buffer1_1/charge_pump1_0/capacitors_1_1/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# cp1_buffer1_2/charge_pump1_0/vdd 3.45f
C692 cp1_buffer1_reverse_1/charge_pump1_reverse_0/capacitor_8_1/capacitor_7_0/buffer_and_gate_0/m1_5444_838# VSUBS 4.07f
C693 cp1_buffer1_reverse_0/charge_pump1_reverse_0/capacitors_1_12/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# cp1_buffer1_2/charge_pump1_0/vdd 13.3f
C694 cp1_buffer1_2/charge_pump1_0/capacitors_1_1/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# cp1_buffer1_2/charge_pump1_0/vdd 3.45f
C695 cp1_buffer1_2/charge_pump1_0/vdd cp1_buffer1_1/charge_pump1_0/capacitors_1_1/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 13.1f
C696 cp1_buffer1_1/charge_pump1_0/capacitors_1_11/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/m1_5444_838# cp1_buffer1_1/charge_pump1_0/capacitors_1_11/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 2.1f
C697 cp1_buffer1_2/charge_pump1_0/vdd cp1_buffer1_0/charge_pump1_0/capacitor_8_1/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 13.3f
C698 cp1_buffer1_2/charge_pump1_0/capacitors_1_1/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/m1_5444_838# cp1_buffer1_2/charge_pump1_0/vdd 8.43f
C699 VSUBS cp1_buffer1_2/charge_pump1_0/capacitors_1_13/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/m1_5444_838# 4.07f
C700 cp1_buffer1_2/charge_pump1_0/m1_12659_300# cp1_buffer1_2/charge_pump1_0/m1_12464_n576# 2.14f
C701 cp1_buffer1_0/charge_pump1_0/capacitors_1_13/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/m1_5444_838# cp1_buffer1_2/charge_pump1_0/vdd 8.43f
C702 cp1_buffer1_reverse_0/charge_pump1_reverse_0/capacitors_1_9/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/m1_5444_838# VSUBS 4.07f
C703 cp1_buffer1_reverse_1/charge_pump1_reverse_0/capacitors_1_11/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# cp1_buffer1_reverse_1/charge_pump1_reverse_0/capacitors_1_11/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/m1_5444_838# 2.1f
C704 cp1_buffer1_0/charge_pump1_0/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/m1_5444_838# cp1_buffer1_2/charge_pump1_0/vdd 8.43f
C705 cp1_buffer1_0/charge_pump1_0/capacitors_1_4/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# cp1_buffer1_2/charge_pump1_0/vdd 13.3f
C706 cp1_buffer1_0/charge_pump1_0/capacitors_1_2/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/m1_5444_838# cp1_buffer1_0/charge_pump1_0/capacitors_1_2/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 2.1f
C707 cp1_buffer1_1/charge_pump1_0/input1 cp1_buffer1_2/charge_pump1_0/vdd 28.3f
C708 cp1_buffer1_2/charge_pump1_0/vdd cp1_buffer1_reverse_1/charge_pump1_reverse_0/nmos_dnw3_0/vs 10.6f
C709 cp1_buffer1_2/charge_pump1_0/input2 VSUBS 10.4f
C710 cp1_buffer1_2/charge_pump1_0/in4 cp1_buffer1_2/charge_pump1_0/capacitors_1_13/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 2.94f
C711 cp1_buffer1_reverse_0/charge_pump1_reverse_0/capacitors_1_7/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/m1_5444_838# VSUBS 4.07f
C712 cp1_buffer1_reverse_0/charge_pump1_reverse_0/capacitors_1_0/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# cp1_buffer1_2/charge_pump1_0/vdd 3.45f
C713 VSUBS cp1_buffer1_1/charge_pump1_0/capacitors_1_3/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/m1_5444_838# 4.07f
C714 cp1_buffer1_reverse_1/charge_pump1_reverse_0/capacitors_1_6/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/m1_5444_838# cp1_buffer1_2/charge_pump1_0/vdd 8.44f
C715 cp1_buffer1_2/charge_pump1_0/in4 cp1_buffer1_reverse_1/charge_pump1_reverse_0/capacitors_1_12/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 2.94f
C716 cp1_buffer1_reverse_0/charge_pump1_reverse_0/capacitor_8_1/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# cp1_buffer1_2/charge_pump1_0/vdd 13.3f
C717 cp1_buffer1_2/charge_pump1_0/capacitors_1_6/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# VSUBS 6.15f
C718 cp1_buffer1_2/charge_pump1_0/capacitors_1_8/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# VSUBS 6.15f
C719 cp1_buffer1_2/charge_pump1_0/vdd cp1_buffer1_0/charge_pump1_0/capacitors_1_8/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# 3.49f
C720 cp1_buffer1_2/charge_pump1_0/in5 cp1_buffer1_reverse_1/charge_pump1_reverse_0/capacitors_1_13/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 2.94f
C721 cp1_buffer1_reverse_1/charge_pump1_reverse_0/capacitors_1_6/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# VSUBS 6.15f
C722 cp1_buffer1_0/charge_pump1_0/clock_0/a_2020_n482# cp1_buffer1_2/charge_pump1_0/vdd 2.66f
C723 cp1_buffer1_reverse_1/charge_pump1_reverse_0/capacitors_1_0/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# VSUBS 6.05f
C724 cp1_buffer1_2/charge_pump1_0/vdd cp1_buffer1_2/charge_pump1_0/capacitors_1_3/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 13.3f
C725 cp1_buffer1_reverse_1/charge_pump1_reverse_0/capacitors_1_6/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# cp1_buffer1_2/charge_pump1_0/vdd 3.49f
C726 cp1_buffer1_reverse_1/charge_pump1_reverse_0/capacitors_1_5/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# cp1_buffer1_reverse_1/charge_pump1_reverse_0/capacitors_1_5/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/m1_5444_838# 2.1f
C727 cp1_buffer1_2/charge_pump1_0/capacitors_1_12/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# cp1_buffer1_2/charge_pump1_0/clkb 2.17f
C728 cp1_buffer1_2/charge_pump1_0/in3 cp1_buffer1_2/charge_pump1_0/capacitors_1_3/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 2.94f
C729 cp1_buffer1_2/charge_pump1_0/in5 cp1_buffer1_1/charge_pump1_0/capacitors_1_7/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 2.94f
C730 cp1_buffer1_2/charge_pump1_0/vdd cp1_buffer1_0/charge_pump1_0/input2 28f
C731 cp1_buffer1_2/charge_pump1_0/vdd cp1_buffer1_1/charge_pump1_0/capacitors_1_8/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# 3.49f
C732 cp1_buffer1_reverse_0/charge_pump1_reverse_0/capacitors_1_13/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/m1_5444_838# cp1_buffer1_2/charge_pump1_0/vdd 8.43f
C733 cp1_buffer1_2/charge_pump1_0/in5 cp1_buffer1_1/charge_pump1_0/capacitors_1_12/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 2.94f
C734 cp1_buffer1_reverse_1/charge_pump1_reverse_0/capacitor_8_1/capacitor_7_0/buffer_and_gate_0/in1 cp1_buffer1_2/charge_pump1_0/in1 2.94f
C735 cp1_buffer1_0/charge_pump1_0/capacitors_1_9/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/m1_5444_838# VSUBS 4.07f
C736 cp1_buffer1_reverse_1/charge_pump1_reverse_0/clock_1/clkb cp1_buffer1_reverse_1/charge_pump1_reverse_0/capacitors_1_9/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 2.17f
C737 cp1_buffer1_1/charge_pump1_0/capacitors_1_10/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# cp1_buffer1_1/charge_pump1_0/capacitors_1_10/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/m1_5444_838# 2.1f
C738 cp1_buffer1_2/charge_pump1_0/vdd cp1_buffer1_2/charge_pump1_0/capacitors_1_12/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# 3.48f
C739 cp1_buffer1_2/charge_pump1_0/vdd cp1_buffer1_1/charge_pump1_0/capacitor_8_1/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 13.3f
C740 VSUBS cp1_buffer1_1/charge_pump1_0/input2 10.4f
C741 cp1_buffer1_2/charge_pump1_0/in4 cp1_buffer1_1/charge_pump1_0/capacitors_1_6/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 2.94f
C742 VSUBS cp1_buffer1_2/charge_pump1_0/clkb 27.8f
C743 cp1_buffer1_2/charge_pump1_0/in3 cp1_buffer1_2/charge_pump1_0/vdd 13.8f
C744 cp1_buffer1_reverse_0/charge_pump1_reverse_0/capacitors_1_13/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# VSUBS 6.15f
C745 cp1_buffer1_reverse_1/charge_pump1_reverse_0/clock_1/clk cp1_buffer1_reverse_1/charge_pump1_reverse_0/input2 8.93f
C746 VSUBS cp1_buffer1_0/charge_pump1_0/capacitors_1_3/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/m1_5444_838# 4.07f
C747 cp1_buffer1_reverse_0/charge_pump1_reverse_0/capacitors_1_13/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# cp1_buffer1_2/charge_pump1_0/vdd 3.48f
C748 cp1_buffer1_1/charge_pump1_0/capacitors_1_9/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# cp1_buffer1_2/charge_pump1_0/vdd 3.48f
C749 cp1_buffer1_0/charge_pump1_0/capacitors_1_4/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# cp1_buffer1_2/charge_pump1_0/vdd 3.48f
C750 cp1_buffer1_0/charge_pump1_0/clkb cp1_buffer1_0/charge_pump1_0/capacitors_1_10/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 2.16f
C751 cp1_buffer1_0/charge_pump1_0/input1 VSUBS 9.98f
C752 cp1_buffer1_0/charge_pump1_0/capacitors_1_5/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/m1_5444_838# VSUBS 4.07f
C753 cp1_buffer1_1/charge_pump1_0/clock_0/a_2402_572# cp1_buffer1_2/charge_pump1_0/vdd 2.67f
C754 cp1_buffer1_2/charge_pump1_0/capacitors_1_4/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# cp1_buffer1_2/charge_pump1_0/vdd 3.48f
C755 cp1_buffer1_1/charge_pump1_0/capacitors_1_7/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# cp1_buffer1_1/charge_pump1_0/capacitors_1_7/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/m1_5444_838# 2.1f
C756 cp1_buffer1_0/charge_pump1_0/capacitors_1_10/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/m1_5444_838# VSUBS 4.07f
C757 cp1_buffer1_reverse_1/charge_pump1_reverse_0/capacitors_1_8/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# cp1_buffer1_2/charge_pump1_0/vdd 13.3f
C758 cp1_buffer1_reverse_1/charge_pump1_reverse_0/capacitors_1_11/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 cp1_buffer1_2/charge_pump1_0/in3 2.94f
C759 cp1_buffer1_1/charge_pump1_0/capacitors_1_12/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# cp1_buffer1_2/charge_pump1_0/vdd 13.3f
C760 cp1_buffer1_0/charge_pump1_0/clk cp1_buffer1_0/charge_pump1_0/capacitors_1_2/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 2.17f
C761 cp1_buffer1_2/charge_pump1_0/capacitors_1_2/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# VSUBS 6.15f
C762 cp1_buffer1_reverse_0/charge_pump1_reverse_0/capacitors_1_10/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# cp1_buffer1_2/charge_pump1_0/vdd 13.3f
C763 cp1_buffer1_1/charge_pump1_0/clk cp1_buffer1_1/charge_pump1_0/input1 8.87f
C764 cp1_buffer1_reverse_1/charge_pump1_reverse_0/capacitors_1_5/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/m1_5444_838# VSUBS 4.07f
C765 cp1_buffer1_2/charge_pump1_0/capacitors_1_2/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/m1_5444_838# cp1_buffer1_2/charge_pump1_0/capacitors_1_2/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 2.1f
C766 cp1_buffer1_1/charge_pump1_0/clk cp1_buffer1_reverse_1/charge_pump1_reverse_0/nmos_dnw3_0/vs 2.31f
C767 cp1_buffer1_2/charge_pump1_0/vin cp1_buffer1_2/charge_pump1_0/vdd 10.3f
C768 cp1_buffer1_reverse_1/charge_pump1_reverse_0/input2 VSUBS 9.75f
C769 cp1_buffer1_reverse_0/charge_pump1_reverse_0/capacitors_1_11/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# cp1_buffer1_reverse_0/charge_pump1_reverse_0/capacitors_1_11/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/m1_5444_838# 2.1f
C770 cp1_buffer1_reverse_0/charge_pump1_reverse_0/capacitors_1_1/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# cp1_buffer1_reverse_0/charge_pump1_reverse_0/clock_1/clk 2.18f
C771 cp1_buffer1_2/charge_pump1_0/in1 cp1_buffer1_1/charge_pump1_0/capacitors_1_0/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 2.94f
C772 cp1_buffer1_2/charge_pump1_0/clk VSUBS 31.5f
C773 cp1_buffer1_reverse_1/charge_pump1_reverse_0/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/m1_5444_838# VSUBS 4.07f
C774 cp1_buffer1_2/charge_pump1_0/in8 cp1_buffer1_0/charge_pump1_0/capacitor_8_1/capacitor_7_0/buffer_and_gate_0/in1 2.94f
C775 cp1_buffer1_reverse_0/charge_pump1_reverse_0/clock_1/a_2432_n962# cp1_buffer1_2/charge_pump1_0/vdd 7.04f
C776 cp1_buffer1_reverse_0/charge_pump1_reverse_0/capacitors_1_8/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/m1_5444_838# cp1_buffer1_2/charge_pump1_0/vdd 8.44f
C777 cp1_buffer1_0/charge_pump1_0/capacitors_1_9/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/m1_5444_838# cp1_buffer1_0/charge_pump1_0/capacitors_1_9/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 2.1f
C778 cp1_buffer1_2/charge_pump1_0/capacitors_1_12/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# cp1_buffer1_2/charge_pump1_0/capacitors_1_12/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/m1_5444_838# 2.1f
C779 cp1_buffer1_2/charge_pump1_0/vdd cp1_buffer1_1/charge_pump1_0/capacitors_1_0/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/m1_5444_838# 8.43f
C780 cp1_buffer1_reverse_0/charge_pump1_reverse_0/capacitors_1_5/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# cp1_buffer1_reverse_0/charge_pump1_reverse_0/capacitors_1_5/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/m1_5444_838# 2.1f
C781 VSUBS cp1_buffer1_2/charge_pump1_0/in7 7.02f
C782 cp1_buffer1_2/charge_pump1_0/in1 cp1_buffer1_2/charge_pump1_0/capacitors_1_0/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 2.94f
C783 cp1_buffer1_reverse_0/charge_pump1_reverse_0/capacitors_1_11/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/m1_5444_838# VSUBS 4.08f
C784 cp1_buffer1_1/charge_pump1_0/clk cp1_buffer1_2/charge_pump1_0/vdd 82.2f
C785 cp1_buffer1_2/charge_pump1_0/clk cp1_buffer1_2/charge_pump1_0/g1 8.15f
C786 cp1_buffer1_reverse_0/charge_pump1_reverse_0/capacitors_1_0/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# VSUBS 6.05f
C787 cp1_buffer1_2/charge_pump1_0/capacitors_1_12/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/m1_5444_838# VSUBS 4.07f
C788 cp1_buffer1_reverse_0/charge_pump1_reverse_0/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# cp1_buffer1_2/charge_pump1_0/vdd 3.48f
C789 VSUBS cp1_buffer1_0/charge_pump1_0/capacitors_1_12/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/m1_5444_838# 4.07f
C790 cp1_buffer1_reverse_0/charge_pump1_reverse_0/input1 cp1_buffer1_2/charge_pump1_0/vdd 27.9f
C791 cp1_buffer1_2/charge_pump1_0/capacitors_1_1/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/m1_5444_838# cp1_buffer1_2/charge_pump1_0/capacitors_1_1/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 2.1f
C792 cp1_buffer1_1/charge_pump1_0/capacitors_1_12/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# cp1_buffer1_2/charge_pump1_0/vdd 3.48f
C793 cp1_buffer1_2/charge_pump1_0/capacitor_8_1/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# cp1_buffer1_2/charge_pump1_0/vdd 3.48f
C794 cp1_buffer1_reverse_1/charge_pump1_reverse_0/capacitors_1_7/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/m1_5444_838# cp1_buffer1_2/charge_pump1_0/vdd 8.44f
Xcp1_buffer1_0/charge_pump1_0 cp1_buffer1_0/charge_pump1_0/clk_in cp1_buffer1_0/charge_pump1_0/input1
+ cp1_buffer1_0/charge_pump1_0/input2 cp1_buffer1_2/charge_pump1_0/vdd VSUBS cp1_buffer1_2/charge_pump1_0/in1
+ cp1_buffer1_2/charge_pump1_0/in3 cp1_buffer1_2/charge_pump1_0/in2 cp1_buffer1_2/charge_pump1_0/in4
+ cp1_buffer1_2/charge_pump1_0/in5 cp1_buffer1_2/charge_pump1_0/in6 cp1_buffer1_2/charge_pump1_0/in7
+ cp1_buffer1_2/charge_pump1_0/in8 cp1_buffer1_0/charge_pump1_0/vin cp1_buffer1_0/charge_pump1_0/g1
+ cp1_buffer1_0/charge_pump1_0/g2 cp1_buffer1_0/charge_pump1_0/clk cp1_buffer1_0/charge_pump1_0/clkb
+ charge_pump1
Xcp1_buffer1_1/charge_pump1_0 cp1_buffer1_1/charge_pump1_0/clk_in cp1_buffer1_1/charge_pump1_0/input1
+ cp1_buffer1_1/charge_pump1_0/input2 cp1_buffer1_2/charge_pump1_0/vdd VSUBS cp1_buffer1_2/charge_pump1_0/in1
+ cp1_buffer1_2/charge_pump1_0/in3 cp1_buffer1_2/charge_pump1_0/in2 cp1_buffer1_2/charge_pump1_0/in4
+ cp1_buffer1_2/charge_pump1_0/in5 cp1_buffer1_2/charge_pump1_0/in6 cp1_buffer1_2/charge_pump1_0/in7
+ cp1_buffer1_2/charge_pump1_0/in8 cp1_buffer1_1/charge_pump1_0/vin cp1_buffer1_1/charge_pump1_0/g1
+ cp1_buffer1_1/charge_pump1_0/g2 cp1_buffer1_1/charge_pump1_0/clk cp1_buffer1_1/charge_pump1_0/clkb
+ charge_pump1
Xcp1_buffer1_2/charge_pump1_0 cp1_buffer1_2/charge_pump1_0/clk_in cp1_buffer1_2/charge_pump1_0/input1
+ cp1_buffer1_2/charge_pump1_0/input2 cp1_buffer1_2/charge_pump1_0/vdd VSUBS cp1_buffer1_2/charge_pump1_0/in1
+ cp1_buffer1_2/charge_pump1_0/in3 cp1_buffer1_2/charge_pump1_0/in2 cp1_buffer1_2/charge_pump1_0/in4
+ cp1_buffer1_2/charge_pump1_0/in5 cp1_buffer1_2/charge_pump1_0/in6 cp1_buffer1_2/charge_pump1_0/in7
+ cp1_buffer1_2/charge_pump1_0/in8 cp1_buffer1_2/charge_pump1_0/vin cp1_buffer1_2/charge_pump1_0/g1
+ cp1_buffer1_2/charge_pump1_0/g2 cp1_buffer1_2/charge_pump1_0/clk cp1_buffer1_2/charge_pump1_0/clkb
+ charge_pump1
Xcp1_buffer1_reverse_0/charge_pump1_reverse_0 cp1_buffer1_2/charge_pump1_0/vdd cp1_buffer1_reverse_0/charge_pump1_reverse_0/input1
+ cp1_buffer1_reverse_0/charge_pump1_reverse_0/input2 VSUBS cp1_buffer1_2/charge_pump1_0/in8
+ cp1_buffer1_2/charge_pump1_0/in6 cp1_buffer1_2/charge_pump1_0/in7 cp1_buffer1_2/charge_pump1_0/in5
+ cp1_buffer1_2/charge_pump1_0/in4 cp1_buffer1_2/charge_pump1_0/in3 cp1_buffer1_2/charge_pump1_0/in2
+ cp1_buffer1_2/charge_pump1_0/in1 charge_pump1_reverse
Xcp1_buffer1_reverse_1/charge_pump1_reverse_0 cp1_buffer1_2/charge_pump1_0/vdd cp1_buffer1_reverse_1/charge_pump1_reverse_0/input1
+ cp1_buffer1_reverse_1/charge_pump1_reverse_0/input2 VSUBS cp1_buffer1_2/charge_pump1_0/in8
+ cp1_buffer1_2/charge_pump1_0/in6 cp1_buffer1_2/charge_pump1_0/in7 cp1_buffer1_2/charge_pump1_0/in5
+ cp1_buffer1_2/charge_pump1_0/in4 cp1_buffer1_2/charge_pump1_0/in3 cp1_buffer1_2/charge_pump1_0/in2
+ cp1_buffer1_2/charge_pump1_0/in1 charge_pump1_reverse
C795 cp1_buffer1_reverse_1/charge_pump1_reverse_0/input1 0 22.9f
C796 cp1_buffer1_reverse_1/charge_pump1_reverse_0/input2 0 22.4f
C797 cp1_buffer1_reverse_1/charge_pump1_reverse_0/capacitors_1_12/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C798 cp1_buffer1_reverse_1/charge_pump1_reverse_0/capacitors_1_12/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C799 cp1_buffer1_reverse_1/charge_pump1_reverse_0/capacitors_1_12/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 0 2.66f
C800 cp1_buffer1_reverse_1/charge_pump1_reverse_0/capacitors_1_13/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C801 cp1_buffer1_reverse_1/charge_pump1_reverse_0/capacitors_1_13/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C802 cp1_buffer1_reverse_1/charge_pump1_reverse_0/capacitors_1_13/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 0 2.66f
C803 cp1_buffer1_reverse_1/charge_pump1_reverse_0/capacitors_1_11/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C804 cp1_buffer1_reverse_1/charge_pump1_reverse_0/capacitors_1_11/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C805 cp1_buffer1_reverse_1/charge_pump1_reverse_0/capacitors_1_11/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 0 2.66f
C806 cp1_buffer1_reverse_1/charge_pump1_reverse_0/capacitors_1_10/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C807 cp1_buffer1_reverse_1/charge_pump1_reverse_0/capacitors_1_10/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C808 cp1_buffer1_reverse_1/charge_pump1_reverse_0/capacitors_1_10/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 0 2.66f
C809 cp1_buffer1_reverse_1/charge_pump1_reverse_0/m1_4341_n519# 0 3.86f
C810 cp1_buffer1_reverse_1/charge_pump1_reverse_0/m1_12659_300# 0 2.73f
C811 cp1_buffer1_2/charge_pump1_0/vin 0 13.3f
C812 cp1_buffer1_reverse_1/charge_pump1_reverse_0/capacitors_1_9/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C813 cp1_buffer1_reverse_1/charge_pump1_reverse_0/capacitors_1_9/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C814 cp1_buffer1_reverse_1/charge_pump1_reverse_0/capacitors_1_9/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 0 2.66f
C815 cp1_buffer1_reverse_1/charge_pump1_reverse_0/capacitors_1_8/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C816 cp1_buffer1_reverse_1/charge_pump1_reverse_0/capacitors_1_8/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C817 cp1_buffer1_reverse_1/charge_pump1_reverse_0/capacitors_1_8/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 0 2.66f
C818 cp1_buffer1_reverse_1/charge_pump1_reverse_0/capacitors_1_7/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C819 cp1_buffer1_reverse_1/charge_pump1_reverse_0/capacitors_1_7/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C820 cp1_buffer1_reverse_1/charge_pump1_reverse_0/capacitors_1_7/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 0 2.66f
C821 cp1_buffer1_2/charge_pump1_0/in4 0 7.84f
C822 cp1_buffer1_reverse_1/charge_pump1_reverse_0/capacitors_1_6/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C823 cp1_buffer1_reverse_1/charge_pump1_reverse_0/capacitors_1_6/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C824 cp1_buffer1_reverse_1/charge_pump1_reverse_0/capacitors_1_6/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 0 2.66f
C825 cp1_buffer1_reverse_1/charge_pump1_reverse_0/capacitors_1_5/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C826 cp1_buffer1_reverse_1/charge_pump1_reverse_0/capacitors_1_5/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C827 cp1_buffer1_reverse_1/charge_pump1_reverse_0/capacitors_1_5/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 0 2.66f
C828 cp1_buffer1_reverse_1/charge_pump1_reverse_0/capacitors_1_4/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C829 cp1_buffer1_reverse_1/charge_pump1_reverse_0/capacitors_1_4/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C830 cp1_buffer1_reverse_1/charge_pump1_reverse_0/capacitors_1_4/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 0 2.66f
C831 cp1_buffer1_reverse_1/charge_pump1_reverse_0/capacitors_1_3/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C832 cp1_buffer1_reverse_1/charge_pump1_reverse_0/capacitors_1_3/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C833 cp1_buffer1_reverse_1/charge_pump1_reverse_0/capacitors_1_3/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 0 2.66f
C834 cp1_buffer1_2/charge_pump1_0/in6 0 7.75f
C835 cp1_buffer1_reverse_1/charge_pump1_reverse_0/capacitors_1_2/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C836 cp1_buffer1_reverse_1/charge_pump1_reverse_0/capacitors_1_2/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C837 cp1_buffer1_reverse_1/charge_pump1_reverse_0/capacitors_1_2/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 0 2.66f
C838 cp1_buffer1_reverse_1/charge_pump1_reverse_0/capacitors_1_1/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C839 cp1_buffer1_reverse_1/charge_pump1_reverse_0/capacitors_1_1/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C840 cp1_buffer1_reverse_1/charge_pump1_reverse_0/capacitors_1_1/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 0 2.66f
C841 cp1_buffer1_reverse_1/charge_pump1_reverse_0/capacitors_1_0/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C842 cp1_buffer1_reverse_1/charge_pump1_reverse_0/capacitors_1_0/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C843 cp1_buffer1_reverse_1/charge_pump1_reverse_0/capacitors_1_0/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 0 2.66f
C844 cp1_buffer1_2/charge_pump1_0/in8 0 8.1f
C845 cp1_buffer1_reverse_1/charge_pump1_reverse_0/capacitor_8_1/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C846 cp1_buffer1_reverse_1/charge_pump1_reverse_0/clock_1/clk 0 88.1f
C847 cp1_buffer1_reverse_1/charge_pump1_reverse_0/capacitor_8_1/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C848 cp1_buffer1_reverse_1/charge_pump1_reverse_0/capacitor_8_1/capacitor_7_0/buffer_and_gate_0/in1 0 2.66f
C849 cp1_buffer1_reverse_1/charge_pump1_reverse_0/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C850 cp1_buffer1_reverse_1/charge_pump1_reverse_0/clock_1/clkb 0 96.8f
C851 cp1_buffer1_reverse_1/charge_pump1_reverse_0/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C852 cp1_buffer1_reverse_1/charge_pump1_reverse_0/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 0 2.66f
C853 cp1_buffer1_reverse_1/charge_pump1_reverse_0/clock_1/a_2432_n962# 0 8.68f
C854 cp1_buffer1_reverse_1/charge_pump1_reverse_0/clock_1/a_2020_n482# 0 2.57f
C855 cp1_buffer1_reverse_1/charge_pump1_reverse_0/clock_1/a_344_102# 0 2.81f **FLOATING
C856 cp1_buffer1_reverse_1/charge_pump1_reverse_0/clock_1/a_2402_572# 0 2.17f
C857 cp1_buffer1_reverse_1/charge_pump1_reverse_0/clock_1/a_344_n986# 0 2.38f **FLOATING
C858 cp1_buffer1_reverse_1/charge_pump1_reverse_0/clock_1/a_3246_118# 0 6.83f
C859 cp1_buffer1_reverse_1/charge_pump1_reverse_0/nmos_dnw3_0/clkb 0 2.01f
C860 cp1_buffer1_reverse_1/charge_pump1_reverse_0/clock_1/clk_in 0 13.9f
C861 cp1_buffer1_reverse_0/charge_pump1_reverse_0/input1 0 22.9f
C862 cp1_buffer1_reverse_0/charge_pump1_reverse_0/input2 0 22.4f
C863 cp1_buffer1_reverse_0/charge_pump1_reverse_0/capacitors_1_12/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C864 cp1_buffer1_reverse_0/charge_pump1_reverse_0/capacitors_1_12/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C865 cp1_buffer1_reverse_0/charge_pump1_reverse_0/capacitors_1_12/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 0 2.66f
C866 cp1_buffer1_reverse_0/charge_pump1_reverse_0/capacitors_1_13/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C867 cp1_buffer1_reverse_0/charge_pump1_reverse_0/capacitors_1_13/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C868 cp1_buffer1_reverse_0/charge_pump1_reverse_0/capacitors_1_13/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 0 2.66f
C869 cp1_buffer1_reverse_0/charge_pump1_reverse_0/capacitors_1_11/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C870 cp1_buffer1_reverse_0/charge_pump1_reverse_0/capacitors_1_11/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C871 cp1_buffer1_reverse_0/charge_pump1_reverse_0/capacitors_1_11/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 0 2.66f
C872 cp1_buffer1_reverse_0/charge_pump1_reverse_0/capacitors_1_10/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C873 cp1_buffer1_reverse_0/charge_pump1_reverse_0/capacitors_1_10/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C874 cp1_buffer1_reverse_0/charge_pump1_reverse_0/capacitors_1_10/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 0 2.66f
C875 cp1_buffer1_reverse_0/charge_pump1_reverse_0/m1_4341_n519# 0 3.86f
C876 cp1_buffer1_reverse_0/charge_pump1_reverse_0/m1_12659_300# 0 2.73f
C877 cp1_buffer1_1/charge_pump1_0/vin 0 13.2f
C878 cp1_buffer1_reverse_0/charge_pump1_reverse_0/capacitors_1_9/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C879 cp1_buffer1_reverse_0/charge_pump1_reverse_0/capacitors_1_9/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C880 cp1_buffer1_reverse_0/charge_pump1_reverse_0/capacitors_1_9/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 0 2.66f
C881 cp1_buffer1_2/charge_pump1_0/in2 0 7.73f
C882 cp1_buffer1_reverse_0/charge_pump1_reverse_0/capacitors_1_8/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C883 cp1_buffer1_reverse_0/charge_pump1_reverse_0/capacitors_1_8/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C884 cp1_buffer1_reverse_0/charge_pump1_reverse_0/capacitors_1_8/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 0 2.66f
C885 cp1_buffer1_reverse_0/charge_pump1_reverse_0/capacitors_1_7/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C886 cp1_buffer1_reverse_0/charge_pump1_reverse_0/capacitors_1_7/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C887 cp1_buffer1_reverse_0/charge_pump1_reverse_0/capacitors_1_7/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 0 2.66f
C888 cp1_buffer1_reverse_0/charge_pump1_reverse_0/capacitors_1_6/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C889 cp1_buffer1_reverse_0/charge_pump1_reverse_0/capacitors_1_6/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C890 cp1_buffer1_reverse_0/charge_pump1_reverse_0/capacitors_1_6/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 0 2.66f
C891 cp1_buffer1_2/charge_pump1_0/in5 0 7.82f
C892 cp1_buffer1_reverse_0/charge_pump1_reverse_0/capacitors_1_5/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C893 cp1_buffer1_reverse_0/charge_pump1_reverse_0/capacitors_1_5/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C894 cp1_buffer1_reverse_0/charge_pump1_reverse_0/capacitors_1_5/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 0 2.66f
C895 cp1_buffer1_reverse_0/charge_pump1_reverse_0/capacitors_1_4/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C896 cp1_buffer1_reverse_0/charge_pump1_reverse_0/capacitors_1_4/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C897 cp1_buffer1_reverse_0/charge_pump1_reverse_0/capacitors_1_4/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 0 2.66f
C898 cp1_buffer1_reverse_0/charge_pump1_reverse_0/capacitors_1_3/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C899 cp1_buffer1_reverse_0/charge_pump1_reverse_0/capacitors_1_3/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C900 cp1_buffer1_reverse_0/charge_pump1_reverse_0/capacitors_1_3/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 0 2.66f
C901 cp1_buffer1_reverse_0/charge_pump1_reverse_0/capacitors_1_2/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C902 cp1_buffer1_reverse_0/charge_pump1_reverse_0/capacitors_1_2/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C903 cp1_buffer1_reverse_0/charge_pump1_reverse_0/capacitors_1_2/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 0 2.66f
C904 cp1_buffer1_reverse_0/charge_pump1_reverse_0/capacitors_1_1/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C905 cp1_buffer1_reverse_0/charge_pump1_reverse_0/capacitors_1_1/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C906 cp1_buffer1_reverse_0/charge_pump1_reverse_0/capacitors_1_1/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 0 2.66f
C907 cp1_buffer1_reverse_0/charge_pump1_reverse_0/capacitors_1_0/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C908 cp1_buffer1_reverse_0/charge_pump1_reverse_0/capacitors_1_0/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C909 cp1_buffer1_reverse_0/charge_pump1_reverse_0/capacitors_1_0/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 0 2.66f
C910 cp1_buffer1_reverse_0/charge_pump1_reverse_0/capacitor_8_1/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C911 cp1_buffer1_reverse_0/charge_pump1_reverse_0/clock_1/clk 0 88.1f
C912 cp1_buffer1_reverse_0/charge_pump1_reverse_0/capacitor_8_1/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C913 cp1_buffer1_reverse_0/charge_pump1_reverse_0/capacitor_8_1/capacitor_7_0/buffer_and_gate_0/in1 0 2.66f
C914 cp1_buffer1_reverse_0/charge_pump1_reverse_0/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C915 cp1_buffer1_reverse_0/charge_pump1_reverse_0/clock_1/clkb 0 96.8f
C916 cp1_buffer1_reverse_0/charge_pump1_reverse_0/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C917 cp1_buffer1_reverse_0/charge_pump1_reverse_0/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 0 2.66f
C918 cp1_buffer1_reverse_0/charge_pump1_reverse_0/clock_1/a_2432_n962# 0 8.68f
C919 cp1_buffer1_reverse_0/charge_pump1_reverse_0/clock_1/a_2020_n482# 0 2.57f
C920 cp1_buffer1_reverse_0/charge_pump1_reverse_0/clock_1/a_344_102# 0 2.81f **FLOATING
C921 cp1_buffer1_reverse_0/charge_pump1_reverse_0/clock_1/a_2402_572# 0 2.17f
C922 cp1_buffer1_reverse_0/charge_pump1_reverse_0/clock_1/a_344_n986# 0 2.38f **FLOATING
C923 cp1_buffer1_reverse_0/charge_pump1_reverse_0/clock_1/a_3246_118# 0 6.83f
C924 cp1_buffer1_reverse_0/charge_pump1_reverse_0/nmos_dnw3_0/clkb 0 2.01f
C925 cp1_buffer1_reverse_0/charge_pump1_reverse_0/clock_1/clk_in 0 10.4f
C926 cp1_buffer1_2/charge_pump1_0/input1 0 22.5f
C927 cp1_buffer1_2/charge_pump1_0/input2 0 22.2f
C928 cp1_buffer1_2/charge_pump1_0/capacitors_1_12/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C929 cp1_buffer1_2/charge_pump1_0/capacitors_1_12/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C930 cp1_buffer1_2/charge_pump1_0/capacitors_1_12/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 0 2.66f
C931 cp1_buffer1_2/charge_pump1_0/capacitors_1_13/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C932 cp1_buffer1_2/charge_pump1_0/capacitors_1_13/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C933 cp1_buffer1_2/charge_pump1_0/capacitors_1_13/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 0 2.66f
C934 cp1_buffer1_2/charge_pump1_0/capacitors_1_11/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C935 cp1_buffer1_2/charge_pump1_0/capacitors_1_11/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C936 cp1_buffer1_2/charge_pump1_0/capacitors_1_11/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 0 2.66f
C937 cp1_buffer1_2/charge_pump1_0/capacitors_1_10/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C938 cp1_buffer1_2/charge_pump1_0/capacitors_1_10/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C939 cp1_buffer1_2/charge_pump1_0/capacitors_1_10/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 0 2.66f
C940 cp1_buffer1_2/charge_pump1_0/m1_4341_n519# 0 3.77f
C941 cp1_buffer1_2/charge_pump1_0/m1_12659_300# 0 2.54f
C942 cp1_buffer1_2/charge_pump1_0/m1_12464_n576# 0 4.25f
C943 cp1_buffer1_2/charge_pump1_0/capacitors_1_9/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C944 cp1_buffer1_2/charge_pump1_0/capacitors_1_9/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C945 cp1_buffer1_2/charge_pump1_0/capacitors_1_9/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 0 2.66f
C946 cp1_buffer1_2/charge_pump1_0/capacitors_1_8/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C947 cp1_buffer1_2/charge_pump1_0/capacitors_1_8/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C948 cp1_buffer1_2/charge_pump1_0/capacitors_1_8/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 0 2.66f
C949 cp1_buffer1_2/charge_pump1_0/capacitors_1_7/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C950 cp1_buffer1_2/charge_pump1_0/capacitors_1_7/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C951 cp1_buffer1_2/charge_pump1_0/capacitors_1_7/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 0 2.66f
C952 cp1_buffer1_2/charge_pump1_0/capacitors_1_6/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C953 cp1_buffer1_2/charge_pump1_0/capacitors_1_6/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C954 cp1_buffer1_2/charge_pump1_0/capacitors_1_6/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 0 2.66f
C955 cp1_buffer1_2/charge_pump1_0/capacitors_1_5/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C956 cp1_buffer1_2/charge_pump1_0/capacitors_1_5/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C957 cp1_buffer1_2/charge_pump1_0/capacitors_1_5/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 0 2.66f
C958 cp1_buffer1_2/charge_pump1_0/capacitors_1_4/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C959 cp1_buffer1_2/charge_pump1_0/capacitors_1_4/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C960 cp1_buffer1_2/charge_pump1_0/capacitors_1_4/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 0 2.66f
C961 cp1_buffer1_2/charge_pump1_0/capacitors_1_3/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C962 cp1_buffer1_2/charge_pump1_0/capacitors_1_3/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C963 cp1_buffer1_2/charge_pump1_0/capacitors_1_3/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 0 2.66f
C964 cp1_buffer1_2/charge_pump1_0/capacitors_1_2/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C965 cp1_buffer1_2/charge_pump1_0/capacitors_1_2/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C966 cp1_buffer1_2/charge_pump1_0/capacitors_1_2/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 0 2.66f
C967 cp1_buffer1_2/charge_pump1_0/capacitors_1_1/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C968 cp1_buffer1_2/charge_pump1_0/capacitors_1_1/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C969 cp1_buffer1_2/charge_pump1_0/capacitors_1_1/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 0 2.66f
C970 cp1_buffer1_2/charge_pump1_0/capacitors_1_0/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C971 cp1_buffer1_2/charge_pump1_0/capacitors_1_0/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C972 cp1_buffer1_2/charge_pump1_0/capacitors_1_0/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 0 2.66f
C973 cp1_buffer1_2/charge_pump1_0/capacitor_8_1/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C974 cp1_buffer1_2/charge_pump1_0/clkb 0 86.1f
C975 cp1_buffer1_2/charge_pump1_0/capacitor_8_1/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C976 cp1_buffer1_2/charge_pump1_0/capacitor_8_1/capacitor_7_0/buffer_and_gate_0/in1 0 2.66f
C977 cp1_buffer1_2/charge_pump1_0/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C978 cp1_buffer1_2/charge_pump1_0/clk 0 85.2f
C979 cp1_buffer1_2/charge_pump1_0/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C980 cp1_buffer1_2/charge_pump1_0/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 0 2.66f
C981 cp1_buffer1_2/charge_pump1_0/clock_0/a_2432_n962# 0 8.68f
C982 cp1_buffer1_2/charge_pump1_0/clock_0/a_2020_n482# 0 2.57f
C983 cp1_buffer1_2/charge_pump1_0/clock_0/a_344_102# 0 2.81f **FLOATING
C984 cp1_buffer1_2/charge_pump1_0/clock_0/a_2402_572# 0 2.17f
C985 cp1_buffer1_2/charge_pump1_0/clock_0/a_344_n986# 0 2.38f **FLOATING
C986 cp1_buffer1_2/charge_pump1_0/clk_in 0 11.3f
C987 cp1_buffer1_2/charge_pump1_0/clock_0/a_3246_118# 0 6.83f
C988 cp1_buffer1_2/charge_pump1_0/g2 0 2.34f
C989 cp1_buffer1_1/charge_pump1_0/input1 0 22.5f
C990 cp1_buffer1_1/charge_pump1_0/input2 0 22.2f
C991 cp1_buffer1_1/charge_pump1_0/capacitors_1_12/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C992 cp1_buffer1_1/charge_pump1_0/capacitors_1_12/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C993 cp1_buffer1_1/charge_pump1_0/capacitors_1_12/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 0 2.66f
C994 cp1_buffer1_1/charge_pump1_0/capacitors_1_13/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C995 cp1_buffer1_1/charge_pump1_0/capacitors_1_13/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C996 cp1_buffer1_1/charge_pump1_0/capacitors_1_13/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 0 2.66f
C997 cp1_buffer1_1/charge_pump1_0/capacitors_1_11/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C998 cp1_buffer1_1/charge_pump1_0/capacitors_1_11/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C999 cp1_buffer1_1/charge_pump1_0/capacitors_1_11/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 0 2.66f
C1000 cp1_buffer1_1/charge_pump1_0/capacitors_1_10/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C1001 cp1_buffer1_1/charge_pump1_0/capacitors_1_10/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C1002 cp1_buffer1_1/charge_pump1_0/capacitors_1_10/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 0 2.66f
C1003 cp1_buffer1_1/charge_pump1_0/m1_4341_n519# 0 3.77f
C1004 cp1_buffer1_1/charge_pump1_0/m1_12659_300# 0 2.54f
C1005 cp1_buffer1_reverse_1/charge_pump1_reverse_0/nmos_dnw3_0/vs 0 14.9f
C1006 cp1_buffer1_1/charge_pump1_0/capacitors_1_9/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C1007 cp1_buffer1_1/charge_pump1_0/capacitors_1_9/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C1008 cp1_buffer1_1/charge_pump1_0/capacitors_1_9/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 0 2.66f
C1009 cp1_buffer1_2/charge_pump1_0/in7 0 7.68f
C1010 cp1_buffer1_1/charge_pump1_0/capacitors_1_8/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C1011 cp1_buffer1_1/charge_pump1_0/capacitors_1_8/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C1012 cp1_buffer1_1/charge_pump1_0/capacitors_1_8/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 0 2.66f
C1013 cp1_buffer1_1/charge_pump1_0/capacitors_1_7/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C1014 cp1_buffer1_1/charge_pump1_0/capacitors_1_7/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C1015 cp1_buffer1_1/charge_pump1_0/capacitors_1_7/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 0 2.66f
C1016 cp1_buffer1_1/charge_pump1_0/capacitors_1_6/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C1017 cp1_buffer1_1/charge_pump1_0/capacitors_1_6/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C1018 cp1_buffer1_1/charge_pump1_0/capacitors_1_6/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 0 2.66f
C1019 cp1_buffer1_1/charge_pump1_0/capacitors_1_5/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C1020 cp1_buffer1_1/charge_pump1_0/capacitors_1_5/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C1021 cp1_buffer1_1/charge_pump1_0/capacitors_1_5/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 0 2.66f
C1022 cp1_buffer1_1/charge_pump1_0/capacitors_1_4/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C1023 cp1_buffer1_1/charge_pump1_0/capacitors_1_4/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C1024 cp1_buffer1_1/charge_pump1_0/capacitors_1_4/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 0 2.66f
C1025 cp1_buffer1_1/charge_pump1_0/capacitors_1_3/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C1026 cp1_buffer1_1/charge_pump1_0/capacitors_1_3/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C1027 cp1_buffer1_1/charge_pump1_0/capacitors_1_3/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 0 2.66f
C1028 cp1_buffer1_2/charge_pump1_0/in3 0 7.71f
C1029 cp1_buffer1_1/charge_pump1_0/capacitors_1_2/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C1030 cp1_buffer1_1/charge_pump1_0/capacitors_1_2/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C1031 cp1_buffer1_1/charge_pump1_0/capacitors_1_2/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 0 2.66f
C1032 cp1_buffer1_1/charge_pump1_0/capacitors_1_1/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C1033 cp1_buffer1_1/charge_pump1_0/capacitors_1_1/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C1034 cp1_buffer1_1/charge_pump1_0/capacitors_1_1/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 0 2.66f
C1035 cp1_buffer1_1/charge_pump1_0/capacitors_1_0/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C1036 cp1_buffer1_1/charge_pump1_0/capacitors_1_0/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C1037 cp1_buffer1_1/charge_pump1_0/capacitors_1_0/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 0 2.66f
C1038 cp1_buffer1_2/charge_pump1_0/in1 0 7.43f
C1039 cp1_buffer1_1/charge_pump1_0/capacitor_8_1/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C1040 cp1_buffer1_1/charge_pump1_0/clkb 0 86.1f
C1041 cp1_buffer1_1/charge_pump1_0/capacitor_8_1/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C1042 cp1_buffer1_1/charge_pump1_0/capacitor_8_1/capacitor_7_0/buffer_and_gate_0/in1 0 2.66f
C1043 cp1_buffer1_1/charge_pump1_0/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C1044 cp1_buffer1_1/charge_pump1_0/clk 0 85.2f
C1045 cp1_buffer1_1/charge_pump1_0/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C1046 cp1_buffer1_1/charge_pump1_0/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 0 2.66f
C1047 cp1_buffer1_1/charge_pump1_0/clock_0/a_2432_n962# 0 8.68f
C1048 cp1_buffer1_1/charge_pump1_0/clock_0/a_2020_n482# 0 2.57f
C1049 cp1_buffer1_1/charge_pump1_0/clock_0/a_344_102# 0 2.81f **FLOATING
C1050 cp1_buffer1_1/charge_pump1_0/clock_0/a_2402_572# 0 2.17f
C1051 cp1_buffer1_1/charge_pump1_0/clock_0/a_344_n986# 0 2.38f **FLOATING
C1052 cp1_buffer1_1/charge_pump1_0/clk_in 0 8.68f
C1053 cp1_buffer1_1/charge_pump1_0/clock_0/a_3246_118# 0 6.83f
C1054 cp1_buffer1_1/charge_pump1_0/g2 0 2.34f
C1055 cp1_buffer1_0/m2_6586_52# 0 3.99f **FLOATING
C1056 cp1_buffer1_0/charge_pump1_0/vin 0 10.4f
C1057 cp1_buffer1_0/charge_pump1_0/input1 0 22.5f
C1058 cp1_buffer1_0/charge_pump1_0/input2 0 22.2f
C1059 cp1_buffer1_0/charge_pump1_0/capacitors_1_12/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C1060 cp1_buffer1_0/charge_pump1_0/capacitors_1_12/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C1061 cp1_buffer1_0/charge_pump1_0/capacitors_1_12/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 0 2.66f
C1062 cp1_buffer1_0/charge_pump1_0/capacitors_1_13/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C1063 cp1_buffer1_0/charge_pump1_0/capacitors_1_13/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C1064 cp1_buffer1_0/charge_pump1_0/capacitors_1_13/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 0 2.66f
C1065 cp1_buffer1_0/charge_pump1_0/capacitors_1_11/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C1066 cp1_buffer1_0/charge_pump1_0/capacitors_1_11/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C1067 cp1_buffer1_0/charge_pump1_0/capacitors_1_11/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 0 2.66f
C1068 cp1_buffer1_0/charge_pump1_0/capacitors_1_10/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C1069 cp1_buffer1_0/charge_pump1_0/capacitors_1_10/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C1070 cp1_buffer1_0/charge_pump1_0/capacitors_1_10/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 0 2.66f
C1071 cp1_buffer1_0/charge_pump1_0/m1_4341_n519# 0 3.77f
C1072 cp1_buffer1_0/charge_pump1_0/m1_12659_300# 0 2.54f
C1073 cp1_buffer1_reverse_0/charge_pump1_reverse_0/nmos_dnw3_0/vs 0 14.6f
C1074 cp1_buffer1_0/charge_pump1_0/capacitors_1_9/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C1075 cp1_buffer1_0/charge_pump1_0/capacitors_1_9/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C1076 cp1_buffer1_0/charge_pump1_0/capacitors_1_9/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 0 2.66f
C1077 cp1_buffer1_0/charge_pump1_0/capacitors_1_8/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C1078 cp1_buffer1_0/charge_pump1_0/capacitors_1_8/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C1079 cp1_buffer1_0/charge_pump1_0/capacitors_1_8/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 0 2.66f
C1080 cp1_buffer1_0/charge_pump1_0/capacitors_1_7/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C1081 cp1_buffer1_0/charge_pump1_0/capacitors_1_7/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C1082 cp1_buffer1_0/charge_pump1_0/capacitors_1_7/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 0 2.66f
C1083 cp1_buffer1_0/charge_pump1_0/capacitors_1_6/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C1084 cp1_buffer1_0/charge_pump1_0/capacitors_1_6/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C1085 cp1_buffer1_0/charge_pump1_0/capacitors_1_6/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 0 2.66f
C1086 cp1_buffer1_0/charge_pump1_0/capacitors_1_5/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C1087 cp1_buffer1_0/charge_pump1_0/capacitors_1_5/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C1088 cp1_buffer1_0/charge_pump1_0/capacitors_1_5/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 0 2.66f
C1089 cp1_buffer1_0/charge_pump1_0/capacitors_1_4/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C1090 cp1_buffer1_0/charge_pump1_0/capacitors_1_4/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C1091 cp1_buffer1_0/charge_pump1_0/capacitors_1_4/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 0 2.66f
C1092 cp1_buffer1_0/charge_pump1_0/capacitors_1_3/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C1093 cp1_buffer1_0/charge_pump1_0/capacitors_1_3/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C1094 cp1_buffer1_0/charge_pump1_0/capacitors_1_3/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 0 2.66f
C1095 cp1_buffer1_0/charge_pump1_0/capacitors_1_2/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C1096 cp1_buffer1_0/charge_pump1_0/capacitors_1_2/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C1097 cp1_buffer1_0/charge_pump1_0/capacitors_1_2/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 0 2.66f
C1098 cp1_buffer1_0/charge_pump1_0/capacitors_1_1/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C1099 cp1_buffer1_0/charge_pump1_0/capacitors_1_1/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C1100 cp1_buffer1_0/charge_pump1_0/capacitors_1_1/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 0 2.66f
C1101 cp1_buffer1_0/charge_pump1_0/capacitors_1_0/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C1102 cp1_buffer1_0/charge_pump1_0/capacitors_1_0/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C1103 cp1_buffer1_0/charge_pump1_0/capacitors_1_0/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 0 2.66f
C1104 cp1_buffer1_0/charge_pump1_0/capacitor_8_1/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C1105 cp1_buffer1_0/charge_pump1_0/clkb 0 86.1f
C1106 cp1_buffer1_0/charge_pump1_0/capacitor_8_1/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C1107 cp1_buffer1_0/charge_pump1_0/capacitor_8_1/capacitor_7_0/buffer_and_gate_0/in1 0 2.66f
C1108 VSUBS 0 0.331p
C1109 cp1_buffer1_0/charge_pump1_0/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C1110 cp1_buffer1_0/charge_pump1_0/clk 0 85.2f
C1111 cp1_buffer1_0/charge_pump1_0/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C1112 cp1_buffer1_2/charge_pump1_0/vdd 0 2.35p
C1113 cp1_buffer1_0/charge_pump1_0/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 0 2.66f
C1114 cp1_buffer1_0/charge_pump1_0/clock_0/a_2432_n962# 0 8.68f
C1115 cp1_buffer1_0/charge_pump1_0/clock_0/a_2020_n482# 0 2.57f
C1116 cp1_buffer1_0/charge_pump1_0/clock_0/a_344_102# 0 2.81f **FLOATING
C1117 cp1_buffer1_0/charge_pump1_0/clock_0/a_2402_572# 0 2.17f
C1118 cp1_buffer1_0/charge_pump1_0/clock_0/a_344_n986# 0 2.38f **FLOATING
C1119 cp1_buffer1_0/charge_pump1_0/clk_in 0 11.8f
C1120 cp1_buffer1_0/charge_pump1_0/clock_0/a_3246_118# 0 6.83f
C1121 cp1_buffer1_0/charge_pump1_0/g2 0 2.34f
