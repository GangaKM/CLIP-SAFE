magic
tech sky130A
magscale 1 2
timestamp 1699423590
<< nwell >>
rect -15174 104225 -12341 104240
rect -15174 101448 161454 104225
rect -15174 100934 -12391 101448
rect 2019 101392 161454 101448
rect -15174 -101697 -12341 100934
rect 1288 -9104 1460 -8793
rect 158621 -101697 161454 101392
rect -15174 -104530 161454 -101697
<< pwell >>
rect 868 -8741 1044 -8525
<< psubdiff >>
rect -18299 107180 -15928 107281
rect 162114 107180 164435 107281
rect -18299 106690 164486 107180
rect -18299 95375 -17534 106690
rect -18198 -102496 -17534 95375
rect -16422 105173 -14905 106690
rect 161678 106286 164486 106690
rect 161678 105173 162589 106286
rect -16422 104758 162589 105173
rect -16422 95375 -15928 104758
rect -16422 -102496 -15964 95375
rect -18198 -104714 -18190 -102496
rect -15972 -104714 -15964 -102496
rect 155796 100790 158000 100809
rect -12010 100168 158000 100790
rect -12010 98854 -11462 100168
rect 155156 99062 158000 100168
rect 155156 98854 156220 99062
rect -12010 98586 156220 98854
rect -11927 97402 -9642 98586
rect -11927 -101312 -11479 97402
rect -10146 -101312 -9642 97402
rect 155796 3296 156220 98586
rect 155768 2849 156220 3296
rect 155768 -2591 156186 2849
rect 155768 -2926 156220 -2591
rect 904 -8613 1000 -8587
rect 904 -8683 936 -8613
rect 975 -8683 1000 -8613
rect 904 -8684 939 -8683
rect 973 -8684 1000 -8683
rect 904 -8702 1000 -8684
rect 155796 -99116 156220 -2926
rect -11927 -101589 -9642 -101312
rect 17961 -99652 156220 -99116
rect 157553 -98458 158000 99062
rect 157553 -99652 157985 -98458
rect 17961 -99717 157985 -99652
rect 17961 -100983 18676 -99717
rect 46170 -100983 157985 -99717
rect 17961 -101329 157985 -100983
rect 162114 96471 162589 104758
rect -18198 -104916 -17534 -104714
rect -18349 -106504 -17534 -104916
rect -16422 -104916 -15964 -104714
rect 162110 -104916 162589 96471
rect -16422 -105695 162589 -104916
rect -16422 -106504 -15512 -105695
rect -18349 -107212 -15512 -106504
rect 161071 -106908 162589 -105695
rect 163701 104758 164486 106286
rect 163701 94820 164435 104758
rect 163701 -104916 164344 94820
rect 163701 -106908 164486 -104916
rect 161071 -107212 164486 -106908
rect -18349 -107893 164486 -107212
<< nsubdiff >>
rect -14661 103067 158938 103707
rect -14661 102035 -14169 103067
rect 158791 102035 158938 103067
rect -14661 101691 158938 102035
rect 159086 102674 161151 103903
rect -14611 101101 -12743 101691
rect -14611 95717 -14316 101101
rect -14735 92859 -14316 95717
rect -14611 -101810 -14316 92859
rect -14647 -103373 -14316 -101810
rect -13136 -101810 -12743 101101
rect 1321 -8876 1415 -8850
rect 1321 -9018 1347 -8876
rect 1389 -9018 1415 -8876
rect 1321 -9042 1415 -9018
rect 159086 -101702 159578 102674
rect 160659 -101702 161151 102674
rect 159086 -101810 161151 -101702
rect -13136 -102411 161151 -101810
rect -13136 -103373 -11982 -102411
rect -14647 -103513 -11982 -103373
rect 159874 -103513 161151 -102411
rect -14647 -104003 161151 -103513
rect 159086 -104013 161151 -104003
<< psubdiffcont >>
rect -17534 -102496 -16422 106690
rect -14905 105173 161678 106690
rect -18190 -104714 -15972 -102496
rect -11462 98854 155156 100168
rect -11479 -101312 -10146 97402
rect 156220 2849 157553 99062
rect 156186 -2591 157553 2849
rect 936 -8683 975 -8613
rect 939 -8684 973 -8683
rect 156220 -99652 157553 -2591
rect 18676 -100983 46170 -99717
rect -17534 -106504 -16422 -104714
rect -15512 -107212 161071 -105695
rect 162589 -106908 163701 106286
<< nsubdiffcont >>
rect -14169 102035 158791 103067
rect -14316 -103373 -13136 101101
rect 1347 -9018 1389 -8876
rect 159578 -101702 160659 102674
rect -11982 -103513 159874 -102411
<< poly >>
rect 148146 1776 148244 1796
rect 148146 1456 148162 1776
rect 148228 1456 148244 1776
rect 148146 1248 148244 1456
rect 148148 562 148246 1124
rect 148150 238 148248 344
rect 148150 136 148170 238
rect 148230 136 148248 238
rect 148150 110 148248 136
<< polycont >>
rect 148162 1456 148228 1776
rect 148170 136 148230 238
<< locali >>
rect -18299 107180 -15928 107281
rect 162114 107180 164435 107281
rect -18299 106690 164486 107180
rect -18299 95375 -17534 106690
rect -22430 3452 -18535 3469
rect -22430 3207 -18510 3452
rect -22430 2324 -22119 3207
rect -19207 2324 -18510 3207
rect -22430 2075 -18510 2324
rect -18918 -110654 -18510 2075
rect -18198 -102496 -17534 95375
rect -18198 -104714 -18190 -102496
rect -18198 -104916 -17534 -104714
rect -18349 -106504 -17534 -104916
rect -16422 105173 -14905 106690
rect 161678 106286 164486 106690
rect 161678 105173 162589 106286
rect -16422 104758 162589 105173
rect -16422 95375 -15928 104758
rect -14736 103067 160953 103736
rect -14736 102035 -14169 103067
rect 158791 102772 160953 103067
rect 158791 102035 159528 102772
rect -14736 101866 159528 102035
rect -14736 101101 -12705 101866
rect -16422 -102496 -15964 95375
rect -14736 94984 -14316 101101
rect -14735 92859 -14316 94984
rect -15972 -104714 -15964 -102496
rect -14575 -103373 -14316 92859
rect -13136 -102107 -12705 101101
rect -11927 100718 -9642 100756
rect -11927 100168 158008 100718
rect -11927 98854 -11462 100168
rect 155156 99062 158008 100168
rect 155156 98854 156220 99062
rect -11927 98538 156220 98854
rect -11927 97402 -9642 98538
rect -11927 -101312 -11479 97402
rect -10146 -101312 -9642 97402
rect 155793 3296 156220 98538
rect 155768 2849 156220 3296
rect 157553 98538 158008 99062
rect 148148 1776 148248 1794
rect 148148 1456 148162 1776
rect 148228 1456 148248 1776
rect 148148 1440 148248 1456
rect 148150 238 148244 254
rect 148150 136 148170 238
rect 148230 136 148244 238
rect 148150 110 148244 136
rect 155768 -2591 156186 2849
rect 155768 -2926 156220 -2591
rect 909 -8613 997 -8589
rect 909 -8683 936 -8613
rect 909 -8684 939 -8683
rect 975 -8683 997 -8613
rect 973 -8684 997 -8683
rect 578 -8713 786 -8695
rect 909 -8702 997 -8684
rect 578 -8763 622 -8713
rect 756 -8742 786 -8713
rect 1269 -8725 1431 -8714
rect 756 -8743 943 -8742
rect 756 -8763 1102 -8743
rect 1269 -8750 1283 -8725
rect 578 -8779 1102 -8763
rect 1136 -8778 1283 -8750
rect 1414 -8778 1431 -8725
rect 578 -8785 786 -8779
rect 1136 -8784 1431 -8778
rect 1321 -8876 1415 -8850
rect 1321 -9018 1347 -8876
rect 1389 -9018 1415 -8876
rect 1321 -9042 1415 -9018
rect 155793 -99106 156220 -2926
rect 44154 -99133 156220 -99106
rect -11927 -101589 -9642 -101312
rect 17972 -99652 156220 -99133
rect 157553 -99106 157979 98538
rect 157553 -99652 157983 -99106
rect 17972 -99698 157983 -99652
rect 17972 -99717 42624 -99698
rect 17972 -99736 18676 -99717
rect 17972 -100999 18658 -99736
rect 157466 -100999 157983 -99698
rect 17972 -101356 157983 -100999
rect 155793 -101388 157979 -101356
rect 159083 -101702 159528 101866
rect 160708 -101702 160953 102772
rect 162114 96471 162589 104758
rect 159083 -102107 160953 -101702
rect -13136 -102411 160953 -102107
rect -13136 -103373 -11982 -102411
rect -14575 -103513 -11982 -103373
rect 159874 -103513 160953 -102411
rect -14575 -103977 160953 -103513
rect -16422 -104916 -15964 -104714
rect 162110 -104916 162589 96471
rect -16422 -105695 162589 -104916
rect -16422 -106504 -15512 -105695
rect -18349 -107212 -15512 -106504
rect 161071 -106908 162589 -105695
rect 163701 104758 164486 106286
rect 163701 94820 164435 104758
rect 163701 -104916 164344 94820
rect 163701 -106908 164486 -104916
rect 161071 -107212 164486 -106908
rect -18349 -107893 164486 -107212
rect -18918 -110928 -12069 -110654
rect -18918 -111747 -18327 -110928
rect -12516 -111747 -12069 -110928
rect -18918 -111995 -12069 -111747
rect -18918 -112075 -18510 -111995
<< viali >>
rect -22119 2324 -19207 3207
rect -17534 -106504 -16422 106690
rect -14905 105173 161678 106690
rect -14169 102035 158791 103067
rect 159528 102674 160708 102772
rect -14316 -103373 -13136 101101
rect -11462 98854 155156 100168
rect -11479 -101312 -10146 97402
rect 156220 2849 157553 99062
rect 148162 1456 148228 1776
rect 148170 136 148230 238
rect 156186 -2591 157553 2849
rect 939 -8684 973 -8614
rect 622 -8763 756 -8713
rect 1283 -8778 1414 -8725
rect 1347 -9018 1389 -8876
rect 156220 -99652 157553 -2591
rect 42624 -99717 157466 -99698
rect 42624 -99736 46170 -99717
rect 18658 -100983 18676 -99736
rect 18676 -100983 46170 -99736
rect 46170 -100983 157466 -99717
rect 18658 -100999 157466 -100983
rect 159528 -101702 159578 102674
rect 159578 -101702 160659 102674
rect 160659 -101702 160708 102674
rect -11982 -103513 159874 -102411
rect -15512 -107212 161071 -105695
rect 162589 -106908 163701 106286
rect -18327 -111747 -12516 -110928
<< metal1 >>
rect -18299 107180 -15928 107281
rect 162114 107180 164435 107281
rect -18299 106690 164486 107180
rect -18299 95375 -17534 106690
rect -22408 3207 -18497 3481
rect -22408 2324 -22119 3207
rect -19207 2324 -18497 3207
rect -22408 2088 -18497 2324
rect -18198 -104916 -17534 95375
rect -18349 -106504 -17534 -104916
rect -16422 105173 -14905 106690
rect 161678 106286 164486 106690
rect 161678 105173 162589 106286
rect -16422 104758 162589 105173
rect -16422 95375 -15928 104758
rect -14653 103671 161041 103760
rect -14653 103067 161066 103671
rect -14653 102035 -14169 103067
rect 158791 102772 161066 103067
rect 158791 102035 159528 102772
rect -14653 101808 159528 102035
rect -14646 101101 -12798 101808
rect -14646 96938 -14316 101101
rect -14725 95717 -14316 96938
rect -16422 -104916 -15964 95375
rect -14735 92859 -14316 95717
rect -14646 -103373 -14316 92859
rect -13136 96938 -12798 101101
rect -11927 100718 -9642 100756
rect -11927 100168 158008 100718
rect -11927 98854 -11462 100168
rect 155156 99062 158008 100168
rect 155156 98854 156220 99062
rect -11927 98538 156220 98854
rect -11927 97402 -9642 98538
rect -13136 92863 -12747 96938
rect -13136 -102046 -12798 92863
rect -11927 -101312 -11479 97402
rect -10146 -99709 -9642 97402
rect -3767 48070 651 48072
rect -6574 47862 651 48070
rect -6574 46716 -3222 47862
rect -3782 -2028 -3222 46716
rect -3782 -5352 -3614 -2028
rect -3246 -5352 -3222 -2028
rect -3782 -48482 -3222 -5352
rect -3052 46572 -2492 46574
rect -3052 46544 440 46572
rect -3052 -6518 -2492 46544
rect -3052 -7226 -2964 -6518
rect -2554 -7226 -2492 -6518
rect -3052 -7300 -2492 -7226
rect -2380 44396 -1820 44402
rect -2380 44368 750 44396
rect -2380 44230 -1820 44368
rect -2380 42908 -2286 44230
rect -1922 42908 -1820 44230
rect -3052 -8660 -2492 -8508
rect -3052 -9368 -2964 -8660
rect -2554 -9368 -2492 -8660
rect -3052 -47164 -2492 -9368
rect -2380 -44988 -1820 42908
rect -1702 43308 -1142 43316
rect -1702 43280 804 43308
rect -1702 42834 -1142 43280
rect -1693 41992 -1142 42834
rect -1693 41586 -1588 41992
rect -1702 40534 -1588 41586
rect -1224 40534 -1142 41992
rect -1016 41744 -474 41752
rect -1016 41740 308 41744
rect -1702 -43900 -1142 40534
rect -1034 41716 308 41740
rect -1034 39544 -474 41716
rect -1034 38202 -1026 39544
rect -526 38202 -474 39544
rect -1034 -42336 -474 38202
rect -352 -41762 208 41136
rect 8730 4374 9252 4388
rect 8660 4316 9252 4374
rect 10397 4352 10537 4358
rect 10388 4346 10552 4352
rect 8660 3350 8916 4316
rect 10290 4182 10552 4346
rect 8606 3276 8962 3350
rect 8606 2824 8662 3276
rect 8896 2824 8962 3276
rect 8606 2784 8962 2824
rect 8730 2782 8802 2784
rect 786 1027 948 1055
rect 786 912 811 1027
rect 922 980 948 1027
rect 922 938 1113 980
rect 922 912 948 938
rect 786 887 948 912
rect 10100 875 10226 3496
rect 10388 2256 10552 4182
rect 12492 4212 13874 4296
rect 12492 3792 12636 4212
rect 13752 3792 13874 4212
rect 12492 3768 13874 3792
rect 148142 3818 148242 3900
rect 12492 3714 14926 3768
rect 13344 3706 14926 3714
rect 148142 3732 151160 3818
rect 10966 3633 11060 3636
rect 14726 3633 14812 3636
rect 10965 3620 14819 3633
rect 10965 3599 10982 3620
rect 10966 3224 10982 3599
rect 11052 3612 14819 3620
rect 11052 3599 14738 3612
rect 11052 3224 11060 3599
rect 10966 3212 11060 3224
rect 14726 2858 14738 3599
rect 14798 3599 14819 3612
rect 14798 2858 14812 3599
rect 14726 2846 14812 2858
rect 148142 3528 148252 3732
rect 151036 3528 151160 3732
rect 148142 3436 151160 3528
rect 14236 2774 14682 2792
rect 14236 2720 14936 2774
rect 14236 2396 14298 2720
rect 14596 2710 14936 2720
rect 14596 2396 14682 2710
rect 14236 2318 14682 2396
rect 10346 2186 10626 2256
rect 10346 1902 10408 2186
rect 10572 1902 10626 2186
rect 10346 1848 10626 1902
rect 148142 1798 148242 3436
rect 155793 3296 156220 98538
rect 155768 2849 156220 3296
rect 157553 98538 158008 99062
rect 151204 1946 152196 2020
rect 148142 1776 148244 1798
rect 148142 1456 148162 1776
rect 148228 1456 148244 1776
rect 151204 1770 151268 1946
rect 152032 1770 152196 1946
rect 151204 1725 152196 1770
rect 151208 1574 151548 1725
rect 151674 1567 152013 1725
rect 148142 1438 148244 1456
rect 9640 838 10226 875
rect 10100 836 10226 838
rect 141714 868 143268 950
rect 148100 945 148136 1242
rect 148264 1160 148394 1168
rect 148264 1138 148320 1160
rect 148254 1108 148320 1138
rect 148384 1108 148394 1160
rect 148254 1104 148394 1108
rect 148264 1098 148394 1104
rect 148264 1096 148346 1098
rect 141714 508 141758 868
rect 143186 508 143268 868
rect 147518 905 148136 945
rect 147518 791 147540 905
rect 147666 791 148136 905
rect 147518 754 148136 791
rect 141714 440 143268 508
rect 148100 496 148136 754
rect 141923 -176 142237 440
rect 148259 384 148298 543
rect 148257 345 148437 384
rect 148150 238 148244 254
rect 148150 136 148170 238
rect 148230 136 148244 238
rect 148150 110 148244 136
rect 9349 -242 14172 -236
rect 9349 -264 14792 -242
rect 9349 -294 14078 -264
rect 9151 -335 14078 -294
rect 9349 -382 14078 -335
rect 14758 -382 14792 -264
rect 9349 -394 14792 -382
rect 9349 -402 14172 -394
rect 15072 -490 147551 -176
rect 10943 -2054 15498 -2019
rect 10943 -2386 10986 -2054
rect 11284 -2386 15498 -2054
rect 148398 -2319 148437 345
rect 151372 382 151468 388
rect 151372 308 151384 382
rect 151456 308 151468 382
rect 151372 296 151468 308
rect 153290 366 153432 394
rect 150720 174 151114 214
rect 150720 68 150748 174
rect 151082 68 151114 174
rect 150720 46 151114 68
rect 151950 -83 152126 -74
rect 151950 -90 152127 -83
rect 151950 -158 151964 -90
rect 152116 -158 152127 -90
rect 151950 -170 152127 -158
rect 152073 -690 152127 -170
rect 152790 -782 152940 192
rect 153290 120 153310 366
rect 153414 120 153432 366
rect 153290 100 153432 120
rect 10943 -2429 15498 -2386
rect 10780 -2892 10848 -2874
rect 10780 -3454 10786 -2892
rect 10457 -3484 10786 -3454
rect 10844 -3454 10848 -2892
rect 15088 -3352 15498 -2429
rect 148384 -2336 154888 -2319
rect 148384 -2375 154901 -2336
rect 148384 -2535 154888 -2375
rect 148384 -2736 154896 -2535
rect 148400 -2952 154896 -2736
rect 155768 -2591 156186 2849
rect 155768 -2926 156220 -2591
rect 10844 -3455 14406 -3454
rect 14458 -3455 14538 -3454
rect 10844 -3484 14727 -3455
rect 10457 -3489 14472 -3484
rect 10457 -3764 14406 -3489
rect 1612 -5797 3583 -5471
rect 1612 -7322 1938 -5797
rect 10457 -6583 10767 -3764
rect 12980 -4086 13876 -3948
rect 12980 -4494 13094 -4086
rect 13714 -4314 13876 -4086
rect 14458 -4228 14472 -3489
rect 14524 -3489 14727 -3484
rect 14524 -4228 14538 -3489
rect 14458 -4242 14538 -4228
rect 14466 -4244 14516 -4242
rect 13714 -4392 14856 -4314
rect 13714 -4494 13876 -4392
rect 12980 -4572 13876 -4494
rect 10994 -5486 11342 -5446
rect 10994 -5800 11040 -5486
rect 11300 -5800 11342 -5486
rect 10994 -5834 11342 -5800
rect 9611 -6645 10767 -6583
rect 9611 -6649 10697 -6645
rect 1612 -7388 1634 -7322
rect 1916 -7388 1938 -7322
rect 1612 -7626 1938 -7388
rect 11057 -7675 11091 -5834
rect 390 -8412 496 -8376
rect 390 -8634 408 -8412
rect 472 -8634 496 -8412
rect 1650 -8478 1976 -8178
rect 911 -8517 1976 -8478
rect 390 -8648 496 -8634
rect 909 -8576 1976 -8517
rect 909 -8614 997 -8576
rect 391 -9024 493 -8648
rect 909 -8684 939 -8614
rect 973 -8684 997 -8614
rect 578 -8710 786 -8695
rect 909 -8702 997 -8684
rect 578 -8763 622 -8710
rect 759 -8742 786 -8710
rect 1269 -8725 1432 -8714
rect 1269 -8726 1283 -8725
rect 1414 -8726 1432 -8725
rect 759 -8743 943 -8742
rect 759 -8763 1102 -8743
rect 1269 -8750 1282 -8726
rect 578 -8779 1102 -8763
rect 578 -8785 786 -8779
rect 1136 -8780 1282 -8750
rect 1420 -8750 1432 -8726
rect 1420 -8780 1434 -8750
rect 1136 -8784 1434 -8780
rect 1331 -8876 1409 -8851
rect 1331 -8975 1347 -8876
rect 1329 -9018 1347 -8975
rect 1389 -8975 1409 -8876
rect 1650 -8919 1976 -8576
rect 1389 -9018 1411 -8975
rect 391 -9126 1128 -9024
rect 1329 -9051 1411 -9018
rect 1191 -9111 1411 -9051
rect 1191 -9114 1410 -9111
rect 1650 -9245 2969 -8919
rect 8486 -9204 9846 -9092
rect 11049 -9204 11121 -8826
rect 8486 -9214 11121 -9204
rect 1650 -9617 1976 -9245
rect 497 -9682 1976 -9617
rect 497 -9892 526 -9682
rect 1804 -9892 1976 -9682
rect 8486 -9776 8602 -9214
rect 9778 -9276 11121 -9214
rect 9778 -9776 9846 -9276
rect 8486 -9846 9846 -9776
rect 497 -9943 1976 -9892
rect -1034 -42364 -118 -42336
rect -1034 -42392 -474 -42364
rect -1702 -43916 384 -43900
rect -1698 -43928 384 -43916
rect -2380 -45006 324 -44988
rect -2360 -45016 324 -45006
rect -3052 -47190 184 -47164
rect -2908 -47192 184 -47190
rect -3782 -48692 545 -48482
rect 155793 -99080 156220 -2926
rect 10473 -99429 14022 -99129
rect 10473 -99709 10773 -99429
rect -10146 -100779 10773 -99709
rect 13547 -99754 14022 -99429
rect 17949 -99652 156220 -99080
rect 157553 -99120 157979 98538
rect 157553 -99652 157985 -99120
rect 17949 -99698 157985 -99652
rect 17949 -99709 42624 -99698
rect 15947 -99736 42624 -99709
rect 15947 -99754 18658 -99736
rect 13547 -100779 18658 -99754
rect -10146 -100999 18658 -100779
rect 157466 -100999 157985 -99698
rect -10146 -101081 157985 -100999
rect -10146 -101312 -9642 -101081
rect 9573 -101104 17446 -101081
rect -11927 -101589 -9642 -101312
rect 17949 -101360 157985 -101081
rect 17949 -101379 157979 -101360
rect 155793 -101388 157979 -101379
rect 159224 -101702 159528 101808
rect 160708 -101702 161066 102772
rect 162114 96471 162589 104758
rect 159224 -102046 161066 -101702
rect -13136 -102104 10523 -102046
rect 15947 -102104 161066 -102046
rect -13136 -102411 161066 -102104
rect -13136 -103373 -11982 -102411
rect -14646 -103513 -11982 -103373
rect 159874 -103513 161066 -102411
rect -14646 -103958 161066 -103513
rect -14513 -103963 161066 -103958
rect 159224 -103989 161066 -103963
rect 162110 -104916 162589 96471
rect -16422 -105681 162589 -104916
rect -16422 -105695 10989 -105681
rect 13851 -105695 162589 -105681
rect -16422 -106504 -15512 -105695
rect -18349 -107212 -15512 -106504
rect 161071 -106908 162589 -105695
rect 163701 104758 164486 106286
rect 163701 94820 164435 104758
rect 163701 -104916 164344 94820
rect 163701 -106908 164486 -104916
rect 161071 -107212 164486 -106908
rect -18349 -107252 10989 -107212
rect 13851 -107252 164486 -107212
rect -18349 -107893 164486 -107252
rect -18198 -108095 -15964 -107893
rect -18798 -110928 -12069 -110654
rect -18798 -111747 -18327 -110928
rect -12516 -111747 -12069 -110928
rect -18798 -111995 -12069 -111747
<< via1 >>
rect -22119 2324 -19207 3207
rect -3614 -5352 -3246 -2028
rect -2964 -7226 -2554 -6518
rect -2286 42908 -1922 44230
rect -2964 -9368 -2554 -8660
rect -1588 40534 -1224 41992
rect -1026 38202 -526 39544
rect 8662 2824 8896 3276
rect 811 912 922 1027
rect 12636 3792 13752 4212
rect 10982 3224 11052 3620
rect 14738 2858 14798 3612
rect 148252 3528 151036 3732
rect 14298 2396 14596 2720
rect 10408 1902 10572 2186
rect 151268 1770 152032 1946
rect 148320 1108 148384 1160
rect 141758 508 143186 868
rect 147540 791 147666 905
rect 148170 136 148230 238
rect 14078 -382 14758 -264
rect 10986 -2386 11284 -2054
rect 151384 308 151456 382
rect 150748 68 151082 174
rect 151964 -158 152116 -90
rect 153310 120 153414 366
rect 10786 -3484 10844 -2892
rect 13094 -4494 13714 -4086
rect 14472 -4228 14524 -3484
rect 11040 -5800 11300 -5486
rect 1634 -7388 1916 -7322
rect 408 -8634 472 -8412
rect 622 -8713 759 -8710
rect 622 -8763 756 -8713
rect 756 -8763 759 -8713
rect 1282 -8778 1283 -8726
rect 1283 -8778 1414 -8726
rect 1414 -8778 1420 -8726
rect 1282 -8780 1420 -8778
rect 526 -9892 1804 -9682
rect 8602 -9776 9778 -9214
rect 10773 -100779 13547 -99429
rect 159607 1871 160669 3056
rect 10989 -105695 13851 -105681
rect 10989 -107212 13851 -105695
rect 10989 -107252 13851 -107212
rect -18327 -111747 -12516 -110928
<< metal2 >>
rect 133308 87497 148018 87509
rect 133308 87428 148020 87497
rect 133308 87269 166338 87428
rect 146558 79019 166338 87269
rect -8551 44230 -1816 44386
rect -8551 42908 -2286 44230
rect -1922 42908 -1816 44230
rect -8551 42824 -1816 42908
rect -8468 41992 -1150 42074
rect -8468 40534 -1588 41992
rect -1224 40534 -1150 41992
rect -8468 40388 -1150 40534
rect -8260 39544 -494 39628
rect -8260 38202 -1026 39544
rect -526 38202 -494 39544
rect -8260 38108 -494 38202
rect -4264 4744 890 7690
rect 8568 6950 11198 7294
rect 8568 5410 8960 6950
rect 10878 5410 11198 6950
rect 8568 5070 11198 5410
rect -22408 3207 -18497 3481
rect -22408 2324 -22119 3207
rect -19207 2324 -18497 3207
rect -22408 2088 -18497 2324
rect -2626 3266 -1628 4744
rect 10674 3980 11034 5070
rect 12520 4212 13874 4286
rect 10668 3636 11056 3980
rect 12520 3792 12636 4212
rect 13752 3792 13874 4212
rect 12520 3712 13874 3792
rect 148146 3732 151160 3818
rect 10668 3620 11060 3636
rect -2626 2398 -2468 3266
rect -1848 2398 -1628 3266
rect 8606 3276 8962 3350
rect 8606 2824 8662 3276
rect 8896 2824 8962 3276
rect 8606 2784 8962 2824
rect 10668 3224 10982 3620
rect 11052 3224 11060 3620
rect 10668 3212 11060 3224
rect 14726 3612 14812 3636
rect -2626 2132 -1628 2398
rect 10346 2186 10626 2256
rect 10346 1902 10408 2186
rect 10572 1902 10626 2186
rect 10346 1848 10626 1902
rect -5184 -680 674 1248
rect 786 1027 948 1055
rect 786 912 811 1027
rect 922 912 948 1027
rect 786 887 948 912
rect 1274 258 1688 260
rect 1156 234 1688 258
rect 1156 126 1198 234
rect 1600 126 1688 234
rect 1156 110 1688 126
rect 1156 108 1348 110
rect 1170 56 1630 58
rect 1156 34 1630 56
rect 1156 -54 1222 34
rect 1596 -54 1630 34
rect 1156 -94 1630 -54
rect -5108 -906 -4096 -680
rect 10668 -806 11056 3212
rect 14726 2858 14738 3612
rect 14798 2858 14812 3612
rect 148146 3528 148252 3732
rect 151036 3528 151160 3732
rect 148146 3436 151160 3528
rect 15833 3272 16533 3315
rect 15833 3184 15888 3272
rect 16384 3184 16533 3272
rect 15833 3149 16533 3184
rect 159058 3056 161125 3278
rect 148400 2983 148817 3023
rect 14726 2846 14812 2858
rect 14236 2720 14682 2792
rect 14236 2396 14298 2720
rect 14596 2396 14682 2720
rect 148370 2667 154640 2983
rect 148370 2566 154648 2667
rect 14236 2318 14682 2396
rect 148378 2250 154648 2566
rect 148383 1168 148425 2250
rect 151204 2019 152196 2020
rect 159058 2019 159607 3056
rect 151203 1946 159607 2019
rect 151203 1770 151268 1946
rect 152032 1871 159607 1946
rect 160669 2019 161125 3056
rect 160669 1871 161171 2019
rect 152032 1770 161171 1871
rect 151203 1680 161171 1770
rect 148312 1160 148425 1168
rect 148312 1138 148320 1160
rect 148254 1108 148320 1138
rect 148384 1108 148425 1160
rect 148254 1104 148425 1108
rect 148312 1098 148425 1104
rect 148383 1097 148425 1098
rect 141714 868 143268 950
rect 141714 508 141758 868
rect 143186 508 143268 868
rect 147518 905 147705 945
rect 147518 791 147540 905
rect 147666 791 147705 905
rect 147518 754 147705 791
rect 141714 440 143268 508
rect 142442 156 142662 440
rect 151372 382 151468 390
rect 151372 308 151384 382
rect 151456 308 151468 382
rect 148148 238 148244 304
rect 12778 -64 147436 156
rect 148148 136 148170 238
rect 148230 142 148244 238
rect 150720 174 151114 214
rect 148230 136 148414 142
rect 148148 46 148414 136
rect 150720 68 150748 174
rect 151082 68 151114 174
rect 150720 46 151114 68
rect 151372 -74 151468 308
rect 153288 366 153436 396
rect 153288 120 153310 366
rect 153414 120 153436 366
rect 151372 -90 152128 -74
rect 151372 -158 151964 -90
rect 152116 -158 152128 -90
rect 151372 -170 152128 -158
rect 14046 -244 14792 -242
rect 153288 -244 153436 120
rect 14046 -264 153436 -244
rect 14046 -382 14078 -264
rect 14758 -382 153436 -264
rect 14046 -392 153436 -382
rect 14046 -394 14792 -392
rect 9786 -894 11056 -806
rect 12788 -808 150818 -588
rect -5108 -1554 -4990 -906
rect -4196 -1554 -4096 -906
rect -5108 -1672 -4096 -1554
rect -3754 -2028 -3176 -1728
rect -3754 -4654 -3614 -2028
rect -3766 -4766 -3614 -4654
rect -3778 -4966 -3614 -4766
rect -3754 -5352 -3614 -4966
rect -3246 -4654 -3176 -2028
rect 1510 -2972 2938 -2926
rect 1510 -3340 1606 -2972
rect 2902 -3340 2938 -2972
rect 1510 -3396 2938 -3340
rect 8528 -2976 9800 -2932
rect 8528 -3338 8576 -2976
rect 9764 -3338 9800 -2976
rect 8528 -3380 9800 -3338
rect -3246 -4966 9188 -4654
rect -3246 -5352 -3176 -4966
rect -3754 -5514 -3176 -5352
rect 8948 -5872 9188 -4966
rect 8948 -5920 9192 -5872
rect 8948 -5922 8982 -5920
rect 8948 -6094 8977 -5922
rect 8948 -6096 8982 -6094
rect 9160 -6096 9192 -5920
rect 8948 -6142 9192 -6096
rect 8948 -6150 9188 -6142
rect -3052 -6518 -2502 -6446
rect -3052 -7126 -2964 -6518
rect -3053 -7204 -2964 -7126
rect -3052 -7226 -2964 -7204
rect -2554 -7126 -2502 -6518
rect 10091 -6750 10344 -894
rect 150598 -1836 150818 -808
rect 152818 -1836 153038 -1276
rect 10943 -2054 11353 -2019
rect 10943 -2386 10986 -2054
rect 11284 -2386 11353 -2054
rect 150598 -2056 153038 -1836
rect 10943 -2429 11353 -2386
rect 10780 -2892 10848 -2874
rect 10780 -3484 10786 -2892
rect 10844 -3484 10848 -2892
rect 10780 -3494 10848 -3484
rect 14458 -3484 14538 -3454
rect 12980 -4086 13876 -3948
rect 12980 -4494 13094 -4086
rect 13714 -4494 13876 -4086
rect 14458 -4228 14472 -3484
rect 14524 -4211 14538 -3484
rect 15850 -3792 16226 -3762
rect 15850 -3920 15898 -3792
rect 16176 -3920 16226 -3792
rect 15850 -3950 16226 -3920
rect 14524 -4228 14710 -4211
rect 14458 -4239 14710 -4228
rect 14458 -4242 14538 -4239
rect 14466 -4244 14516 -4242
rect 12980 -4572 13876 -4494
rect 10994 -5486 11342 -5446
rect 10994 -5800 11040 -5486
rect 11300 -5800 11342 -5486
rect 10994 -5834 11342 -5800
rect -2554 -7204 2318 -7126
rect -2554 -7226 -2502 -7204
rect -3052 -7308 -2502 -7226
rect 71 -7322 1941 -7303
rect 71 -7388 1634 -7322
rect 1916 -7388 1941 -7322
rect 71 -7410 1941 -7388
rect 71 -8378 178 -7410
rect 71 -8412 498 -8378
rect 71 -8485 408 -8412
rect -3048 -8660 -2498 -8572
rect 391 -8634 408 -8485
rect 472 -8634 498 -8412
rect 391 -8653 498 -8634
rect -3048 -8696 -2964 -8660
rect -3052 -8788 -2964 -8696
rect -3048 -9368 -2964 -8788
rect -2554 -8696 -2498 -8660
rect -2554 -8710 788 -8696
rect -2554 -8763 622 -8710
rect 759 -8763 788 -8710
rect 1270 -8726 1432 -8714
rect 1270 -8750 1282 -8726
rect -2554 -8788 788 -8763
rect 1206 -8780 1282 -8750
rect 1420 -8750 1432 -8726
rect 1420 -8780 2246 -8750
rect 1206 -8784 2246 -8780
rect -2554 -9368 -2498 -8788
rect -3048 -9434 -2498 -9368
rect 8486 -9214 9846 -9092
rect 420 -9682 1968 -9586
rect 420 -9704 526 -9682
rect -4326 -9892 526 -9704
rect 1804 -9892 1968 -9682
rect 8486 -9776 8602 -9214
rect 9778 -9776 9846 -9214
rect 8486 -9846 9846 -9776
rect -4326 -9940 1968 -9892
rect -4326 -12110 1058 -9940
rect 161022 -80316 166580 -79794
rect 147308 -87889 166580 -80316
rect 132474 -88070 166580 -87889
rect 132474 -88129 148006 -88070
rect 147370 -88143 148000 -88129
rect 10473 -99429 14022 -99129
rect 10473 -100779 10773 -99429
rect 13547 -100779 14022 -99429
rect 10473 -101079 14022 -100779
rect 10583 -105681 14586 -104896
rect 10583 -107252 10989 -105681
rect 13851 -107252 14586 -105681
rect 10583 -107936 14586 -107252
rect -18798 -110928 -12069 -110654
rect -18798 -111747 -18327 -110928
rect -12516 -111747 -12069 -110928
rect -18798 -111995 -12069 -111747
<< via2 >>
rect 8960 5410 10878 6950
rect -22119 2324 -19207 3207
rect 12636 3792 13752 4212
rect -2468 2398 -1848 3266
rect 8662 2824 8896 3276
rect 10408 1902 10572 2186
rect 811 912 922 1027
rect 1198 126 1600 234
rect 1222 -54 1596 34
rect 148252 3528 151036 3732
rect 15888 3184 16384 3272
rect 14298 2396 14596 2720
rect 151268 1770 152032 1946
rect 141758 508 143186 868
rect 147540 791 147666 905
rect 150748 68 151082 174
rect -4990 -1554 -4196 -906
rect 1606 -3340 2902 -2972
rect 8576 -3338 9764 -2976
rect 8982 -5922 9160 -5920
rect 8977 -6094 9160 -5922
rect 8982 -6096 9160 -6094
rect 10986 -2386 11284 -2054
rect 10786 -3484 10844 -2892
rect 13094 -4494 13714 -4086
rect 15898 -3920 16176 -3792
rect 11040 -5800 11300 -5486
rect 526 -9892 1804 -9682
rect 8602 -9776 9778 -9214
rect 10773 -100779 13547 -99429
rect 10989 -107252 13851 -105681
rect -18327 -111747 -12516 -110928
<< metal3 >>
rect -8526 6950 11258 7274
rect -8526 5410 8960 6950
rect 10878 5410 11258 6950
rect -8526 5070 11258 5410
rect -22408 3207 -18497 3481
rect -5176 3446 -2824 3456
rect -5176 3444 -824 3446
rect -22408 2324 -22119 3207
rect -19207 2324 -18497 3207
rect -22408 2088 -18497 2324
rect -5178 3266 -824 3444
rect -5178 3222 -2468 3266
rect -5178 2274 -4942 3222
rect -3104 2398 -2468 3222
rect -1848 2398 -824 3266
rect 8606 3276 8962 3350
rect 8606 2824 8662 3276
rect 8896 2824 8962 3276
rect 8606 2784 8962 2824
rect -3104 2276 -824 2398
rect -3104 2274 706 2276
rect -5178 1392 706 2274
rect 10346 2186 10626 2256
rect 10346 1902 10408 2186
rect 10572 1902 10626 2186
rect 10346 1848 10626 1902
rect -4218 1384 -824 1392
rect -6585 1027 948 1054
rect -6585 912 811 1027
rect 922 912 948 1027
rect -6585 888 948 912
rect 8294 802 8906 876
rect -6570 522 1696 591
rect -6582 392 1696 454
rect -6582 329 1699 392
rect -6584 258 1138 264
rect 1274 260 1390 264
rect 1274 258 1688 260
rect -6584 234 1688 258
rect -6584 136 1198 234
rect 1070 126 1198 136
rect 1600 126 1688 234
rect 1070 110 1688 126
rect 1088 48 1222 50
rect 1088 36 1630 48
rect -6575 34 1630 36
rect -6575 -54 1222 34
rect 1596 -54 1630 34
rect -6575 -94 1630 -54
rect -6575 -98 1222 -94
rect 10564 -375 10828 -374
rect 9549 -450 10851 -375
rect -5104 -906 780 -784
rect -5104 -1554 -4990 -906
rect -4196 -1554 780 -906
rect -5104 -1668 780 -1554
rect -104 -2878 780 -1668
rect -104 -2896 2032 -2878
rect -104 -2972 3252 -2896
rect -104 -3340 1606 -2972
rect 2902 -3340 3252 -2972
rect -104 -3454 3252 -3340
rect 8492 -2976 9900 -2888
rect 8492 -3338 8576 -2976
rect 9764 -3338 9900 -2976
rect 8492 -3448 9900 -3338
rect 10564 -2892 10851 -450
rect 10943 -2054 11353 -2019
rect 10943 -2386 10986 -2054
rect 11284 -2386 11353 -2054
rect 10943 -2429 11353 -2386
rect 10564 -3484 10786 -2892
rect 10844 -3484 10851 -2892
rect 8949 -5872 9188 -5868
rect 8948 -5920 9192 -5872
rect 8948 -5922 8982 -5920
rect 8948 -6094 8977 -5922
rect 8948 -6096 8982 -6094
rect 9160 -6096 9192 -5920
rect 8948 -6142 9192 -6096
rect 8949 -6143 9188 -6142
rect 8486 -9214 9846 -9092
rect 420 -9682 1968 -9586
rect 420 -9892 526 -9682
rect 1804 -9892 1968 -9682
rect 8486 -9776 8602 -9214
rect 9778 -9776 9846 -9214
rect 8486 -9846 9846 -9776
rect 420 -9940 1968 -9892
rect 10564 -10166 10851 -3484
rect 10994 -5486 11342 -5446
rect 10994 -5800 11040 -5486
rect 11300 -5800 11342 -5486
rect 10994 -5834 11342 -5800
rect -11674 -11775 10851 -10166
rect -11674 -11810 10710 -11775
rect 9785 -30482 11338 -30481
rect 11530 -30482 12425 30261
rect 12520 4212 13874 4286
rect 12520 3792 12636 4212
rect 13752 3792 13874 4212
rect 12520 3712 13874 3792
rect 15833 3272 16452 3314
rect 15833 3184 15888 3272
rect 16384 3184 16452 3272
rect 15833 3149 16452 3184
rect 14236 2720 14682 2792
rect 14236 2396 14298 2720
rect 14596 2396 14682 2720
rect 14236 2318 14682 2396
rect 141714 868 143268 950
rect 141714 508 141758 868
rect 143186 508 143268 868
rect 141714 440 143268 508
rect 147523 905 147705 6789
rect 148146 3732 151160 3818
rect 148146 3528 148252 3732
rect 151036 3528 151160 3732
rect 148146 3436 151160 3528
rect 151204 1946 152196 2020
rect 151204 1770 151268 1946
rect 152032 1770 152196 1946
rect 151204 1725 152196 1770
rect 147523 791 147540 905
rect 147666 791 147705 905
rect 142650 232 143030 440
rect 147523 232 147705 791
rect 142650 174 151159 232
rect 142650 68 150748 174
rect 151082 68 151159 174
rect 142650 50 151159 68
rect 142650 -140 143030 50
rect 15062 -520 147620 -140
rect 142551 -1206 144558 -1108
rect 151336 -1204 151438 -1014
rect 149920 -1206 151438 -1204
rect 142264 -1210 151438 -1206
rect 142264 -1410 142634 -1210
rect 144396 -1310 151438 -1210
rect 144396 -1410 151378 -1310
rect 142264 -1502 151378 -1410
rect 15850 -3792 16226 -3762
rect 15850 -3824 15898 -3792
rect 15755 -3885 15898 -3824
rect 15850 -3920 15898 -3885
rect 16176 -3920 16226 -3792
rect 12980 -4086 13876 -3948
rect 15850 -3950 16226 -3920
rect 12980 -4494 13094 -4086
rect 13714 -4494 13876 -4086
rect 12980 -4572 13876 -4494
rect 9785 -31539 12425 -30482
rect 9785 -33235 10843 -31539
rect -12084 -95510 10770 -87288
rect 10473 -99429 14022 -99129
rect 10473 -100779 10773 -99429
rect 13547 -100779 14022 -99429
rect 10473 -101079 14022 -100779
rect 10583 -105681 14586 -104896
rect 10583 -107252 10989 -105681
rect 13851 -107252 14586 -105681
rect 10583 -107936 14586 -107252
rect -18798 -110928 -12069 -110654
rect -18798 -111747 -18327 -110928
rect -12516 -111747 -12069 -110928
rect -18798 -111995 -12069 -111747
<< via3 >>
rect -22119 2324 -19207 3207
rect -4942 2274 -3104 3222
rect -2468 2398 -1848 3266
rect 8662 2824 8896 3276
rect 10408 1902 10572 2186
rect -4990 -1554 -4196 -906
rect 8576 -3338 9764 -2976
rect 10986 -2386 11284 -2054
rect 8977 -6094 9155 -5922
rect 526 -9892 1804 -9682
rect 8602 -9776 9778 -9214
rect 11040 -5800 11300 -5486
rect 12636 3792 13752 4212
rect 14298 2396 14596 2720
rect 141758 508 143186 868
rect 148252 3528 151036 3732
rect 151268 1770 152032 1946
rect 142634 -1410 144396 -1210
rect 13094 -4494 13714 -4086
rect 10773 -100779 13547 -99429
rect 10989 -107252 13851 -105681
rect -18327 -111747 -12516 -110928
<< metal4 >>
rect -42087 103024 17476 108254
rect -42087 98072 17648 103024
rect 16921 94385 17619 98072
rect -4264 4744 890 7690
rect -22408 3207 -18497 3481
rect -22408 2324 -22119 3207
rect -19207 2324 -18497 3207
rect -22408 2088 -18497 2324
rect -5176 3222 -2824 3456
rect -5176 2274 -4942 3222
rect -3104 2274 -2824 3222
rect -5176 2076 -2824 2274
rect -2626 3266 -1628 4744
rect 12492 4212 13874 4296
rect 12492 3792 12636 4212
rect 13752 3792 13874 4212
rect 12492 3714 13874 3792
rect -2626 2398 -2468 3266
rect -1848 2398 -1628 3266
rect 8606 3278 8962 3350
rect 8606 2824 8654 3278
rect 8910 2824 8962 3278
rect 8606 2784 8962 2824
rect 14276 2788 14684 2794
rect -2626 2132 -1628 2398
rect 14238 2720 14684 2788
rect 14238 2396 14298 2720
rect 14596 2396 14684 2720
rect 14238 2252 14684 2396
rect 9102 2186 14684 2252
rect 9102 1902 10408 2186
rect 10572 1902 14684 2186
rect 9102 1844 14684 1902
rect -5190 -682 1060 1212
rect 10930 128 11338 1844
rect 141714 868 143268 950
rect 141714 508 141758 868
rect 143186 508 143268 868
rect 141714 440 143268 508
rect 140356 128 141376 178
rect -5108 -906 -4096 -682
rect -5108 -1554 -4990 -906
rect -4196 -1554 -4096 -906
rect -5108 -1672 -4096 -1554
rect 10930 -866 141618 128
rect 10930 -2019 11338 -866
rect 140268 -870 141376 -866
rect 140268 -1102 141272 -870
rect 140268 -1210 144598 -1102
rect 140268 -1410 142634 -1210
rect 144396 -1410 144598 -1210
rect 140268 -1492 144598 -1410
rect 10930 -2054 11353 -2019
rect 10930 -2386 10986 -2054
rect 11284 -2386 11353 -2054
rect 10930 -2429 11353 -2386
rect 8492 -2976 9900 -2888
rect -10346 -4062 -4938 -3018
rect 8492 -3338 8576 -2976
rect 9764 -3338 9900 -2976
rect 8492 -3448 9900 -3338
rect 10930 -4062 11338 -2429
rect -10346 -4470 11338 -4062
rect -10346 -4950 -4938 -4470
rect 10930 -5432 11338 -4470
rect 12980 -4086 13876 -3948
rect 12980 -4494 13094 -4086
rect 13714 -4494 13876 -4086
rect 12980 -4572 13876 -4494
rect 8528 -5486 11338 -5432
rect 8528 -5800 11040 -5486
rect 11300 -5800 11338 -5486
rect 8528 -5840 11338 -5800
rect 8946 -5922 9195 -5904
rect 8946 -6094 8977 -5922
rect 9155 -6094 9195 -5922
rect 8946 -6430 9195 -6094
rect 145536 -7134 146104 4496
rect 148146 3732 151152 4574
rect 148146 3528 148252 3732
rect 151036 3528 151152 3732
rect 148146 3436 151152 3528
rect 151204 1946 152196 2020
rect 151204 1770 151268 1946
rect 152032 1770 152196 1946
rect 151204 1725 152196 1770
rect 151204 -700 151550 1725
rect 8486 -9214 9846 -9092
rect 420 -9682 1968 -9586
rect 420 -9704 526 -9682
rect -4326 -9892 526 -9704
rect 1804 -9892 1968 -9682
rect 8486 -9776 8602 -9214
rect 9778 -9776 9846 -9214
rect 8486 -9846 9846 -9776
rect -4326 -9940 1968 -9892
rect -4326 -12110 1058 -9940
rect 10473 -99429 14022 -99129
rect 10473 -100779 10773 -99429
rect 13547 -100779 14022 -99429
rect 10473 -101079 14022 -100779
rect 10583 -105681 14586 -104896
rect 10583 -107252 10989 -105681
rect 13851 -107252 14586 -105681
rect 10583 -107936 14586 -107252
rect -18798 -110928 -12069 -110654
rect -18798 -111747 -18327 -110928
rect -12516 -111747 -12069 -110928
rect -18798 -111995 -12069 -111747
rect -12432 -113425 -6589 -112623
rect -12432 -114424 -11561 -113425
rect -13282 -114761 -11561 -114424
rect -12432 -115281 -11561 -114761
rect -7941 -115281 -6589 -113425
rect -12432 -116014 -6589 -115281
<< via4 >>
rect -22119 2324 -19207 3207
rect -4942 2274 -3104 3222
rect 12636 3792 13752 4212
rect -2468 2398 -1848 3266
rect 8654 3276 8910 3278
rect 8654 2824 8662 3276
rect 8662 2824 8896 3276
rect 8896 2824 8910 3276
rect 141758 508 143186 868
rect 8576 -3338 9764 -2976
rect 13094 -4494 13714 -4086
rect 8602 -9776 9778 -9214
rect 10773 -100779 13547 -99429
rect 10989 -107252 13851 -105681
rect -18327 -111747 -12516 -110928
rect -11561 -115281 -7941 -113425
<< metal5 >>
rect 146169 5724 146682 5849
rect 12502 4212 13877 4293
rect 12502 3792 12636 4212
rect 13752 3792 13877 4212
rect -22408 3463 -18497 3481
rect 12502 3463 13877 3792
rect -22408 3278 13877 3463
rect -22408 3266 8654 3278
rect -22408 3222 -2468 3266
rect -22408 3207 -4942 3222
rect -22408 2324 -22119 3207
rect -19207 2324 -4942 3207
rect -22408 2274 -4942 2324
rect -3104 2398 -2468 3222
rect -1848 2824 8654 3266
rect 8910 2824 13877 3278
rect -1848 2398 13877 2824
rect -3104 2274 13877 2398
rect -22408 2088 13877 2274
rect 8483 -2702 9858 2088
rect 141714 944 143268 950
rect 138862 868 143292 944
rect 138862 508 141758 868
rect 143186 508 143292 868
rect 138862 442 143292 508
rect 13033 82 13831 297
rect 138874 82 140192 442
rect 141714 440 143268 442
rect 13033 -786 141618 82
rect 8480 -2726 9860 -2702
rect 13033 -2726 13831 -786
rect 138874 -852 140192 -786
rect 8458 -2976 13866 -2726
rect 8458 -3338 8576 -2976
rect 9764 -3338 13866 -2976
rect 8458 -3524 13866 -3338
rect 8480 -9214 9860 -3524
rect 12983 -4086 13866 -3524
rect 12983 -4494 13094 -4086
rect 13714 -4494 13866 -4086
rect 12983 -4559 13866 -4494
rect 12983 -4565 13781 -4559
rect 146169 -7895 146759 5724
rect 8480 -9776 8602 -9214
rect 9778 -9776 9860 -9214
rect 8480 -10294 9860 -9776
rect 15603 -98230 16321 -97802
rect -12568 -99429 16452 -98230
rect -12568 -100779 10773 -99429
rect 13547 -100779 16452 -99429
rect -12568 -105681 16452 -100779
rect -12568 -107252 10989 -105681
rect 13851 -107252 16452 -105681
rect -12568 -109101 16452 -107252
rect -12596 -110641 16511 -109101
rect -18778 -110654 16511 -110641
rect -18798 -110928 16511 -110654
rect -18798 -111747 -18327 -110928
rect -12516 -111747 16511 -110928
rect -18798 -111995 16511 -111747
rect -18778 -112016 16511 -111995
rect -12596 -113425 16511 -112016
rect -12596 -115281 -11561 -113425
rect -7941 -115281 16511 -113425
rect -12596 -116321 16511 -115281
use cmfb_pmos  cmfb_pmos_0 ~/layout_files/differential_amplifier
timestamp 1699272401
transform 1 0 148450 0 1 -716
box -158 762 4965 2374
use comparator_final_compact  comparator_final_compact_0 ~/layout_files/differential_amplifier
timestamp 1699409311
transform -1 0 8641 0 1 -7048
box -2532 -2214 8653 1614
use full_stage_compact  full_stage_compact_0 ~/layout_files/differential_amplifier
timestamp 1699256576
transform 1 0 5194 0 1 -2632
box -4134 -770 6100 4979
use reconfigurable_CP  reconfigurable_CP_0
timestamp 1699265676
transform 1 0 16242 0 -1 63194
box -16084 -34774 130792 62844
use reconfigurable_CP  reconfigurable_CP_1
timestamp 1699265676
transform 1 0 15920 0 1 -63814
box -16084 -34774 130792 62844
use reference0_9  reference0_9_0
timestamp 1699232519
transform 0 -1 151950 1 0 -1600
box -66 -1120 1022 620
use reference  reference_0 ~/layout_files/differential_amplifier
timestamp 1699232519
transform 0 1 9900 -1 0 4400
box -32 -858 1956 500
use sky130_fd_pr__cap_mim_m3_1_LJ5JLG  sky130_fd_pr__cap_mim_m3_1_LJ5JLG_0
timestamp 1699146224
transform -1 0 150592 0 -1 7074
box -3186 -3040 3186 3040
use sky130_fd_pr__nfet_01v8_PXJ6TW  sky130_fd_pr__nfet_01v8_PXJ6TW_0
timestamp 1699271609
transform 1 0 148196 0 1 1206
box -108 -126 108 126
use sky130_fd_pr__nfet_01v8_PXJ6TW  sky130_fd_pr__nfet_01v8_PXJ6TW_1
timestamp 1699271609
transform 1 0 148198 0 1 446
box -108 -126 108 126
use sky130_fd_sc_hd__inv_1  sky130_fd_sc_hd__inv_1_0 ~/sky_pdk/sky130/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1693170804
transform -1 0 1266 0 -1 -8521
box -38 -48 314 592
use source_follower_buffer  source_follower_buffer_0
timestamp 1698922888
transform 1 0 14893 0 1 -4323
box -217 -59 950 1017
use source_follower_buffer  source_follower_buffer_1
timestamp 1698922888
transform 1 0 14975 0 -1 3723
box -217 -59 950 1017
<< labels >>
flabel metal5 15603 -105367 15617 -105363 0 FreeSans 4800 90 0 0 digital_gnd
flabel metal4 16921 102321 17619 103019 0 FreeSans 4800 90 0 0 digital_vdd
rlabel metal3 1158 358 1158 358 1 source
flabel space 8228 39660 9060 39802 0 FreeSans 3200 0 0 0 scan_out
flabel space 148376 1942 148438 2082 0 FreeSans 2400 90 0 0 vd1
flabel space 148306 -658 148460 -292 0 FreeSans 2400 90 0 0 vd2
flabel metal4 -30725 98072 -20543 108254 0 FreeSans 16000 0 0 0 digital_vdd_1.8V
flabel space -6158 -95630 2366 -87288 0 FreeSans 16000 0 0 0 clock(internal)_50MHz
flabel metal5 -6522 -108146 -1140 -101858 0 FreeSans 16000 0 0 0 Digital_gnd
flabel metal2 157929 79019 166338 87428 0 FreeSans 16000 0 0 0 vout+
flabel metal2 153340 2296 153890 2902 0 FreeSans 8000 0 0 0 vd1
flabel space 153456 -2960 154006 -2354 0 FreeSans 8000 0 0 0 vd2
flabel space 153424 -88070 161700 -79794 0 FreeSans 16000 0 0 0 vout-
flabel space -6574 46716 -5648 48142 0 FreeSans 8000 0 0 0 clk_external
flabel metal2 -7251 42824 -5689 44386 0 FreeSans 8000 0 0 0 scan_in
flabel metal2 -8468 40388 -6658 42012 0 FreeSans 8000 0 0 0 scan_en
flabel metal2 -8260 38108 -6042 39556 0 FreeSans 8000 0 0 0 reset
flabel space -5816 -100 -5606 34 0 FreeSans 1600 0 0 0 drain1
flabel space -5822 136 -5612 270 0 FreeSans 1600 0 0 0 drain2
rlabel metal3 1220 550 1220 550 1 ib1
rlabel space -5788 314 -5664 458 1 source
flabel space -5792 310 -5656 472 0 FreeSans 1600 0 0 0 source
flabel space -5886 612 -5706 680 0 FreeSans 1600 0 0 0 ib1
flabel space -5812 1068 -5638 1152 0 FreeSans 1600 0 0 0 ib2_1uA
flabel psubdiff -11610 -11898 -9966 -10254 0 FreeSans 8000 0 0 0 v_int-
flabel metal3 -8526 5070 -6322 7274 0 FreeSans 8000 0 0 0 v_int+
flabel space -10456 2110 -8262 3522 0 FreeSans 6400 0 0 0 analog_gnd
flabel metal4 -10346 -4950 -8000 -3018 0 FreeSans 6400 0 0 0 analog_vdd_1.8V
rlabel via1 912 962 912 962 1 ib2
<< end >>
