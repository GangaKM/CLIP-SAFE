* SPICE3 file created from comparator_full_compact.ext - technology: sky130A

.subckt sky130_fd_pr__pfet_01v8_BH9SS5 w_n246_n319# a_n50_n197# a_50_n100# a_n108_n100#
+ VSUBS
X0 a_50_n100# a_n50_n197# a_n108_n100# w_n246_n319# sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
C0 w_n246_n319# a_n50_n197# 0.279f
C1 a_n50_n197# a_n108_n100# 0.0163f
C2 w_n246_n319# a_50_n100# 0.0852f
C3 a_50_n100# a_n108_n100# 0.0906f
C4 w_n246_n319# a_n108_n100# 0.0852f
C5 a_50_n100# a_n50_n197# 0.0163f
C6 a_50_n100# VSUBS 0.0558f
C7 a_n108_n100# VSUBS 0.0558f
C8 a_n50_n197# VSUBS 0.179f
C9 w_n246_n319# VSUBS 1.41f
.ends

.subckt sky130_fd_pr__nfet_01v8_53744R a_n210_n274# a_50_n100# a_n108_n100# a_n50_n188#
X0 a_50_n100# a_n50_n188# a_n108_n100# a_n210_n274# sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
C0 a_n50_n188# a_n108_n100# 0.0163f
C1 a_n108_n100# a_50_n100# 0.0906f
C2 a_n50_n188# a_50_n100# 0.0163f
C3 a_50_n100# a_n210_n274# 0.141f
C4 a_n108_n100# a_n210_n274# 0.141f
C5 a_n50_n188# a_n210_n274# 0.443f
.ends

.subckt inverter m1_176_134# m1_272_214# li_n18_880# VSUBS
Xsky130_fd_pr__pfet_01v8_BH9SS5_0 li_n18_880# m1_176_134# m1_272_214# li_n18_880#
+ VSUBS sky130_fd_pr__pfet_01v8_BH9SS5
Xsky130_fd_pr__nfet_01v8_53744R_0 VSUBS m1_272_214# VSUBS m1_176_134# sky130_fd_pr__nfet_01v8_53744R
C0 li_n18_880# m1_176_134# 0.137f
C1 li_n18_880# m1_272_214# -0.0185f
C2 m1_272_214# m1_176_134# 0.404f
C3 m1_272_214# VSUBS 0.241f
C4 m1_176_134# VSUBS 0.76f
C5 li_n18_880# VSUBS 1.47f
.ends

.subckt sky130_fd_pr__nfet_01v8_PVEW3M a_n210_n274# a_50_n100# a_n108_n100# a_n50_n188#
X0 a_50_n100# a_n50_n188# a_n108_n100# a_n210_n274# sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
C0 a_50_n100# a_n108_n100# 0.0906f
C1 a_n108_n100# a_n50_n188# 0.0163f
C2 a_50_n100# a_n50_n188# 0.0163f
C3 a_50_n100# a_n210_n274# 0.141f
C4 a_n108_n100# a_n210_n274# 0.141f
C5 a_n50_n188# a_n210_n274# 0.443f
.ends

.subckt sky130_fd_pr__pfet_01v8_X3YSY6 w_n246_n319# a_n50_n197# a_50_n100# a_n108_n100#
+ VSUBS
X0 a_50_n100# a_n50_n197# a_n108_n100# w_n246_n319# sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
C0 a_50_n100# w_n246_n319# 0.0852f
C1 a_n108_n100# a_n50_n197# 0.0163f
C2 a_n50_n197# w_n246_n319# 0.279f
C3 a_n108_n100# w_n246_n319# 0.0852f
C4 a_n50_n197# a_50_n100# 0.0163f
C5 a_n108_n100# a_50_n100# 0.0906f
C6 a_50_n100# VSUBS 0.0558f
C7 a_n108_n100# VSUBS 0.0558f
C8 a_n50_n197# VSUBS 0.179f
C9 w_n246_n319# VSUBS 1.41f
.ends

.subckt sky130_fd_pr__pfet_01v8_B5E2Q5 w_n246_n319# a_n50_n197# a_50_n100# a_n108_n100#
+ VSUBS
X0 a_50_n100# a_n50_n197# a_n108_n100# w_n246_n319# sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
C0 a_50_n100# w_n246_n319# 0.0852f
C1 a_n108_n100# a_n50_n197# 0.0163f
C2 a_n50_n197# w_n246_n319# 0.279f
C3 a_n108_n100# w_n246_n319# 0.0852f
C4 a_n50_n197# a_50_n100# 0.0163f
C5 a_n108_n100# a_50_n100# 0.0906f
C6 a_50_n100# VSUBS 0.0558f
C7 a_n108_n100# VSUBS 0.0558f
C8 a_n50_n197# VSUBS 0.179f
C9 w_n246_n319# VSUBS 1.41f
.ends

.subckt comparator_layout m1_1704_1482# m1_1411_1896# m1_2488_2128# li_905_2237# m1_2014_1251#
+ XM33/a_n50_n188# XM34/a_n50_n188# m1_1061_1257# m1_852_1342# VSUBS XM25/a_n50_n188#
+ XM26/a_n50_n188#
XXM34 VSUBS m1_852_1342# m1_2014_1251# XM34/a_n50_n188# sky130_fd_pr__nfet_01v8_PVEW3M
XXM35 VSUBS VSUBS m1_852_1342# m1_2488_2128# sky130_fd_pr__nfet_01v8_PVEW3M
XXM25 VSUBS m1_1061_1257# m1_852_1342# XM25/a_n50_n188# sky130_fd_pr__nfet_01v8_PVEW3M
XXM26 VSUBS m1_1061_1257# m1_852_1342# XM26/a_n50_n188# sky130_fd_pr__nfet_01v8_PVEW3M
XXM27 VSUBS m1_1411_1896# m1_1061_1257# m1_1704_1482# sky130_fd_pr__nfet_01v8_PVEW3M
XXM28 VSUBS m1_1704_1482# m1_2014_1251# m1_1411_1896# sky130_fd_pr__nfet_01v8_PVEW3M
XXM29 li_905_2237# m1_2488_2128# m1_1411_1896# li_905_2237# VSUBS sky130_fd_pr__pfet_01v8_X3YSY6
Xsky130_fd_pr__pfet_01v8_B5E2Q5_0 li_905_2237# m1_2488_2128# m1_2014_1251# m1_1061_1257#
+ VSUBS sky130_fd_pr__pfet_01v8_B5E2Q5
XXM30 li_905_2237# m1_1704_1482# m1_1411_1896# li_905_2237# VSUBS sky130_fd_pr__pfet_01v8_X3YSY6
XXM31 li_905_2237# m1_1411_1896# m1_1704_1482# li_905_2237# VSUBS sky130_fd_pr__pfet_01v8_X3YSY6
XXM32 li_905_2237# m1_2488_2128# m1_1704_1482# li_905_2237# VSUBS sky130_fd_pr__pfet_01v8_X3YSY6
XXM33 VSUBS m1_852_1342# m1_2014_1251# XM33/a_n50_n188# sky130_fd_pr__nfet_01v8_PVEW3M
C0 m1_852_1342# m1_1061_1257# 0.178f
C1 m1_1704_1482# li_905_2237# 0.438f
C2 m1_2488_2128# XM33/a_n50_n188# 0.0212f
C3 m1_1411_1896# XM33/a_n50_n188# 0.0158f
C4 XM26/a_n50_n188# m1_2014_1251# 5.12e-19
C5 XM26/a_n50_n188# XM25/a_n50_n188# 0.0158f
C6 m1_1061_1257# m1_2014_1251# 0.158f
C7 m1_1061_1257# XM25/a_n50_n188# 0.0289f
C8 li_905_2237# XM33/a_n50_n188# 0.00867f
C9 m1_2488_2128# m1_852_1342# 0.288f
C10 m1_1411_1896# m1_852_1342# 0.0265f
C11 m1_1704_1482# XM33/a_n50_n188# 0.0119f
C12 XM26/a_n50_n188# m1_1061_1257# 0.0834f
C13 m1_2488_2128# XM34/a_n50_n188# 0.0244f
C14 m1_852_1342# li_905_2237# 0.0843f
C15 li_905_2237# XM34/a_n50_n188# 0.00553f
C16 m1_852_1342# m1_1704_1482# 0.0464f
C17 m1_2488_2128# m1_2014_1251# 0.208f
C18 m1_1411_1896# m1_2014_1251# 0.128f
C19 m1_1704_1482# XM34/a_n50_n188# 9.68e-19
C20 li_905_2237# m1_2014_1251# 0.0933f
C21 li_905_2237# XM25/a_n50_n188# 0.00558f
C22 m1_2488_2128# XM26/a_n50_n188# 0.0134f
C23 m1_1411_1896# XM26/a_n50_n188# 7.18e-21
C24 m1_2488_2128# m1_1061_1257# 0.618f
C25 m1_1411_1896# m1_1061_1257# 0.105f
C26 m1_852_1342# XM33/a_n50_n188# 0.0284f
C27 m1_1704_1482# m1_2014_1251# 0.0992f
C28 XM26/a_n50_n188# li_905_2237# 0.00553f
C29 li_905_2237# m1_1061_1257# 0.183f
C30 XM33/a_n50_n188# XM34/a_n50_n188# 0.0158f
C31 m1_1704_1482# XM26/a_n50_n188# 0.0158f
C32 m1_1704_1482# m1_1061_1257# 0.626f
C33 XM33/a_n50_n188# m1_2014_1251# 0.0409f
C34 m1_852_1342# XM34/a_n50_n188# 0.0758f
C35 m1_1411_1896# m1_2488_2128# 0.22f
C36 m1_2488_2128# li_905_2237# 0.747f
C37 m1_852_1342# m1_2014_1251# 0.86f
C38 m1_852_1342# XM25/a_n50_n188# 0.0359f
C39 m1_1411_1896# li_905_2237# 0.48f
C40 m1_1061_1257# XM33/a_n50_n188# 0.0104f
C41 m1_2488_2128# m1_1704_1482# 0.313f
C42 m1_2014_1251# XM34/a_n50_n188# 0.0491f
C43 m1_1411_1896# m1_1704_1482# 0.795f
C44 m1_852_1342# XM26/a_n50_n188# 0.0222f
C45 XM33/a_n50_n188# VSUBS 0.478f
C46 m1_1704_1482# VSUBS 0.845f
C47 m1_1411_1896# VSUBS 0.836f
C48 m1_2488_2128# VSUBS 1.37f
C49 li_905_2237# VSUBS 6.29f
C50 m1_2014_1251# VSUBS 0.749f
C51 XM26/a_n50_n188# VSUBS 0.474f
C52 m1_1061_1257# VSUBS 0.739f
C53 m1_852_1342# VSUBS 2.36f
C54 XM25/a_n50_n188# VSUBS 0.478f
C55 XM34/a_n50_n188# VSUBS 0.474f
.ends

.subckt latch_layout m1_724_1961# m1_1878_998# m1_827_1096# m1_1097_1325# m1_430_1104#
+ m1_822_1732# m1_1595_1096# m1_330_1963# m1_1878_1968# li_30_2070# m1_1601_1730#
+ VSUBS
XXM23 VSUBS m1_430_1104# m1_827_1096# m1_1097_1325# sky130_fd_pr__nfet_01v8_PVEW3M
XXM24 VSUBS m1_1595_1096# m1_1097_1325# m1_430_1104# sky130_fd_pr__nfet_01v8_PVEW3M
XXM14 li_30_2070# m1_724_1961# m1_822_1732# li_30_2070# VSUBS sky130_fd_pr__pfet_01v8_X3YSY6
XXM13 li_30_2070# m1_330_1963# m1_430_1104# li_30_2070# VSUBS sky130_fd_pr__pfet_01v8_X3YSY6
XXM15 li_30_2070# m1_1097_1325# m1_430_1104# m1_822_1732# VSUBS sky130_fd_pr__pfet_01v8_X3YSY6
XXM16 li_30_2070# m1_430_1104# m1_1601_1730# m1_1097_1325# VSUBS sky130_fd_pr__pfet_01v8_X3YSY6
XXM17 li_30_2070# m1_1878_1968# li_30_2070# m1_1601_1730# VSUBS sky130_fd_pr__pfet_01v8_X3YSY6
XXM19 VSUBS VSUBS m1_1595_1096# m1_1878_998# sky130_fd_pr__nfet_01v8_PVEW3M
Xsky130_fd_pr__pfet_01v8_X3YSY6_0 li_30_2070# m1_1878_998# li_30_2070# m1_1097_1325#
+ VSUBS sky130_fd_pr__pfet_01v8_X3YSY6
XXM20 VSUBS VSUBS m1_1097_1325# m1_1878_1968# sky130_fd_pr__nfet_01v8_PVEW3M
XXM21 VSUBS m1_430_1104# VSUBS m1_724_1961# sky130_fd_pr__nfet_01v8_PVEW3M
XXM22 VSUBS m1_827_1096# VSUBS m1_330_1963# sky130_fd_pr__nfet_01v8_PVEW3M
C0 m1_822_1732# m1_827_1096# 0.024f
C1 m1_822_1732# m1_330_1963# 0.00173f
C2 li_30_2070# m1_1097_1325# 0.467f
C3 m1_822_1732# m1_430_1104# -0.0453f
C4 m1_1097_1325# m1_1601_1730# 0.0928f
C5 m1_827_1096# m1_330_1963# 8.98e-20
C6 m1_827_1096# m1_430_1104# -0.0404f
C7 m1_822_1732# m1_724_1961# 3e-20
C8 m1_430_1104# m1_1595_1096# 0.134f
C9 li_30_2070# m1_1601_1730# 0.107f
C10 m1_1097_1325# m1_1878_998# 0.0882f
C11 m1_1878_1968# m1_1097_1325# 0.222f
C12 m1_430_1104# m1_330_1963# 0.136f
C13 m1_330_1963# m1_724_1961# 0.225f
C14 m1_430_1104# m1_724_1961# 0.36f
C15 li_30_2070# m1_1878_998# 0.294f
C16 m1_1878_1968# li_30_2070# 0.152f
C17 m1_1878_998# m1_1601_1730# 4.26e-19
C18 m1_1878_1968# m1_1601_1730# 0.00552f
C19 m1_822_1732# m1_1097_1325# 0.117f
C20 m1_1878_1968# m1_1878_998# 0.258f
C21 m1_1097_1325# m1_827_1096# 0.134f
C22 m1_1097_1325# m1_1595_1096# -0.0527f
C23 m1_822_1732# li_30_2070# 0.105f
C24 li_30_2070# m1_827_1096# 0.0114f
C25 m1_1097_1325# m1_330_1963# 0.0496f
C26 m1_1097_1325# m1_430_1104# 1.73f
C27 li_30_2070# m1_1595_1096# 0.0108f
C28 m1_1601_1730# m1_1595_1096# 0.0228f
C29 m1_1097_1325# m1_724_1961# 0.0408f
C30 m1_822_1732# m1_1878_998# 5.25e-20
C31 li_30_2070# m1_330_1963# 0.193f
C32 li_30_2070# m1_430_1104# 0.32f
C33 m1_1601_1730# m1_330_1963# 1.5e-19
C34 m1_1601_1730# m1_430_1104# 0.0908f
C35 li_30_2070# m1_724_1961# 0.149f
C36 m1_1878_998# m1_1595_1096# 0.00175f
C37 m1_1878_1968# m1_1595_1096# 0.00131f

C38 m1_1878_998# m1_330_1963# 0.00409f
C39 m1_1878_1968# m1_330_1963# 5.9e-20
C40 m1_1878_998# m1_430_1104# 0.0556f
C41 m1_1878_1968# m1_430_1104# 0.0418f
C42 m1_1878_998# m1_724_1961# 0.0025f
C43 m1_1878_1968# m1_724_1961# 0.00416f
C44 m1_1878_998# VSUBS 1.37f
C45 m1_724_1961# VSUBS 0.62f
C46 m1_827_1096# VSUBS 0.309f
C47 m1_1878_1968# VSUBS 0.646f
C48 m1_1601_1730# VSUBS 0.0344f
C49 m1_1097_1325# VSUBS 1.37f
C50 m1_430_1104# VSUBS 1.32f
C51 m1_330_1963# VSUBS 1.27f
C52 li_30_2070# VSUBS 7.27f
C53 m1_822_1732# VSUBS 0.0351f
C54 m1_1595_1096# VSUBS 0.307f
.ends

.subckt comparator_full_compact Vdd gnd clk Vc- V+ V- Vc+ Q Q1
Xinverter_0 vo- vo1- Vdd gnd inverter
Xinverter_1 vo+ vo1+ Vdd gnd inverter
Xcomparator_layout_0 vo- vo+ clk Vdd m1_2098_364# V- Vc- m1_950_364# comparator_layout_0/m1_852_1342#
+ gnd Vc+ V+ comparator_layout
Xlatch_layout_0 vo1+ vo+ latch_layout_0/m1_827_1096# Q1 Q latch_layout_0/m1_822_1732#
+ latch_layout_0/m1_1595_1096# vo- vo1- Vdd latch_layout_0/m1_1601_1730# gnd latch_layout
C0 vo1- Vc- 4.21e-22
C1 Q1 Vc- 4.22e-20
C2 V- clk 0.00182f
C3 vo1+ vo1- 2.5f
C4 vo+ comparator_layout_0/m1_852_1342# 0.00803f
C5 Vc- vo- -3.08e-19
C6 Vdd V- 0.00689f
C7 m1_950_364# V+ 0.0192f
C8 vo1+ vo- 1.27f
C9 vo1+ Vc+ 4.71e-20
C10 Q clk 0.00281f
C11 m1_950_364# vo+ 0.015f
C12 vo1- comparator_layout_0/m1_852_1342# 3.78e-19
C13 m1_2098_364# Vc- 0.0391f
C14 Vdd clk 0.092f
C15 Q1 comparator_layout_0/m1_852_1342# 1.2e-20
C16 Vdd Q 0.00821f
C17 vo- comparator_layout_0/m1_852_1342# 0.0425f
C18 Vc+ comparator_layout_0/m1_852_1342# 0.0347f
C19 vo1- m1_950_364# 9.72e-20
C20 Q1 m1_950_364# 3.33e-22
C21 latch_layout_0/m1_822_1732# clk 5.15e-22
C22 V+ vo+ 0.00406f
C23 m1_2098_364# comparator_layout_0/m1_852_1342# 0.00885f
C24 m1_950_364# vo- 0.0311f
C25 Vc- V- 1.98e-19
C26 latch_layout_0/m1_822_1732# Vdd 5.19e-19
C27 m1_950_364# Vc+ 4.93e-20
C28 vo1+ V- 4.71e-22
C29 latch_layout_0/m1_1601_1730# Vdd -0.00136f
C30 vo1- V+ 4.21e-22
C31 m1_950_364# m1_2098_364# 0.00401f
C32 Vc- clk 2.26e-21
C33 vo1+ clk 0.0256f
C34 Vdd Vc- 8.01e-23
C35 V+ vo- 2.51e-19
C36 latch_layout_0/m1_1595_1096# vo+ 0.00298f
C37 vo1+ Q 0.00149f
C38 vo1- vo+ 0.396f
C39 V+ Vc+ 1.6e-19
C40 vo1+ Vdd 0.664f
C41 Q1 vo+ 0.0506f
C42 vo+ vo- 0.859f
C43 vo+ Vc+ 0.00398f
C44 clk comparator_layout_0/m1_852_1342# -1.48e-19
C45 m1_950_364# V- 0.00162f
C46 Q comparator_layout_0/m1_852_1342# 0.00805f
C47 vo1- Q1 0.104f
C48 Vdd comparator_layout_0/m1_852_1342# -0.00185f
C49 m1_2098_364# vo+ 0.0503f
C50 vo1- vo- 0.025f
C51 m1_950_364# clk 6.92e-19
C52 vo1- Vc+ 4.21e-20
C53 m1_950_364# Q 2.03e-19
C54 latch_layout_0/m1_827_1096# vo+ 0.00298f
C55 m1_950_364# Vdd 7.66e-19
C56 Vc+ vo- 0.0268f
C57 vo1+ Vc- 4.71e-22
C58 Q1 m1_2098_364# 1.21e-20
C59 vo+ V- 0.00427f
C60 m1_2098_364# vo- 0.111f
C61 V+ clk -5.78e-21
C62 Vdd V+ 1.11e-22
C63 Vc- comparator_layout_0/m1_852_1342# 0.0236f
C64 vo+ clk 0.155f
C65 vo1+ comparator_layout_0/m1_852_1342# 8.88e-19
C66 vo1- V- 4.21e-22
C67 vo+ Q 0.028f
C68 Vdd vo+ 0.956f
C69 m1_950_364# Vc- 8.32e-19
C70 V- vo- 0.00101f
C71 vo1+ m1_950_364# 5.47e-20
C72 vo1- clk 0.00428f
C73 Q1 clk 2e-19
C74 vo1- Q 0.0217f
C75 vo1- Vdd 0.594f
C76 Q1 Q 0.00302f
C77 latch_layout_0/m1_822_1732# vo+ 0.0162f
C78 Q1 Vdd -0.00217f
C79 m1_2098_364# V- 0.0328f
C80 clk vo- 0.64f
C81 Q vo- 0.00561f
C82 Vdd vo- 1.2f
C83 latch_layout_0/m1_1601_1730# vo+ 0.0117f
C84 m1_950_364# comparator_layout_0/m1_852_1342# -0.0115f
C85 Vdd Vc+ 0.00363f
C86 vo1+ V+ 4.71e-22
C87 m1_2098_364# clk -0.00123f
C88 latch_layout_0/m1_822_1732# vo1- 0.00386f
C89 latch_layout_0/m1_822_1732# Q1 2.84e-32
C90 m1_2098_364# Q 2.54e-19
C91 Vc- vo+ 0.00413f
C92 Vdd m1_2098_364# 0.0148f
C93 vo1- latch_layout_0/m1_1601_1730# 0.00583f
C94 vo1+ vo+ 0.402f
C95 latch_layout_0/m1_827_1096# Vdd 3.12e-22
C96 V+ comparator_layout_0/m1_852_1342# 0.0302f
C97 latch_layout_0/m1_827_1096# gnd 0.214f
C98 vo1- gnd 2.22f
C99 latch_layout_0/m1_1601_1730# gnd 0.0321f
C100 Q1 gnd 0.985f
C101 Q gnd 0.945f
C102 latch_layout_0/m1_822_1732# gnd 0.0326f
C103 latch_layout_0/m1_1595_1096# gnd 0.213f
C104 V- gnd 0.448f
C105 vo- gnd 2.12f
C106 vo+ gnd 3.92f
C107 clk gnd 0.842f
C108 Vdd gnd 14.6f
C109 m1_2098_364# gnd 0.498f
C110 V+ gnd 0.446f
C111 m1_950_364# gnd 0.496f
C112 comparator_layout_0/m1_852_1342# gnd 1.39f
C113 Vc+ gnd 0.434f
C114 Vc- gnd 0.446f
C115 vo1+ gnd 0.951f
.ends

