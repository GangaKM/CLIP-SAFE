magic
tech sky130A
magscale 1 2
timestamp 1698095665
<< nmos >>
rect -399 -42 -369 42
rect -303 -42 -273 42
rect -207 -42 -177 42
rect -111 -42 -81 42
rect -15 -42 15 42
rect 81 -42 111 42
rect 177 -42 207 42
rect 273 -42 303 42
rect 369 -42 399 42
<< ndiff >>
rect -461 30 -399 42
rect -461 -30 -449 30
rect -415 -30 -399 30
rect -461 -42 -399 -30
rect -369 30 -303 42
rect -369 -30 -353 30
rect -319 -30 -303 30
rect -369 -42 -303 -30
rect -273 30 -207 42
rect -273 -30 -257 30
rect -223 -30 -207 30
rect -273 -42 -207 -30
rect -177 30 -111 42
rect -177 -30 -161 30
rect -127 -30 -111 30
rect -177 -42 -111 -30
rect -81 30 -15 42
rect -81 -30 -65 30
rect -31 -30 -15 30
rect -81 -42 -15 -30
rect 15 30 81 42
rect 15 -30 31 30
rect 65 -30 81 30
rect 15 -42 81 -30
rect 111 30 177 42
rect 111 -30 127 30
rect 161 -30 177 30
rect 111 -42 177 -30
rect 207 30 273 42
rect 207 -30 223 30
rect 257 -30 273 30
rect 207 -42 273 -30
rect 303 30 369 42
rect 303 -30 319 30
rect 353 -30 369 30
rect 303 -42 369 -30
rect 399 30 461 42
rect 399 -30 415 30
rect 449 -30 461 30
rect 399 -42 461 -30
<< ndiffc >>
rect -449 -30 -415 30
rect -353 -30 -319 30
rect -257 -30 -223 30
rect -161 -30 -127 30
rect -65 -30 -31 30
rect 31 -30 65 30
rect 127 -30 161 30
rect 223 -30 257 30
rect 319 -30 353 30
rect 415 -30 449 30
<< poly >>
rect -321 114 -255 130
rect -321 80 -305 114
rect -271 80 -255 114
rect -399 42 -369 68
rect -321 64 -255 80
rect -129 114 -63 130
rect -129 80 -113 114
rect -79 80 -63 114
rect -303 42 -273 64
rect -207 42 -177 68
rect -129 64 -63 80
rect 63 114 129 130
rect 63 80 79 114
rect 113 80 129 114
rect -111 42 -81 64
rect -15 42 15 68
rect 63 64 129 80
rect 255 114 321 130
rect 255 80 271 114
rect 305 80 321 114
rect 81 42 111 64
rect 177 42 207 68
rect 255 64 321 80
rect 273 42 303 64
rect 369 42 399 68
rect -399 -64 -369 -42
rect -417 -80 -351 -64
rect -303 -68 -273 -42
rect -207 -64 -177 -42
rect -417 -114 -401 -80
rect -367 -114 -351 -80
rect -417 -130 -351 -114
rect -225 -80 -159 -64
rect -111 -68 -81 -42
rect -15 -64 15 -42
rect -225 -114 -209 -80
rect -175 -114 -159 -80
rect -225 -130 -159 -114
rect -33 -80 33 -64
rect 81 -68 111 -42
rect 177 -64 207 -42
rect -33 -114 -17 -80
rect 17 -114 33 -80
rect -33 -130 33 -114
rect 159 -80 225 -64
rect 273 -68 303 -42
rect 369 -64 399 -42
rect 159 -114 175 -80
rect 209 -114 225 -80
rect 159 -130 225 -114
rect 351 -80 417 -64
rect 351 -114 367 -80
rect 401 -114 417 -80
rect 351 -130 417 -114
<< polycont >>
rect -305 80 -271 114
rect -113 80 -79 114
rect 79 80 113 114
rect 271 80 305 114
rect -401 -114 -367 -80
rect -209 -114 -175 -80
rect -17 -114 17 -80
rect 175 -114 209 -80
rect 367 -114 401 -80
<< locali >>
rect -321 80 -305 114
rect -271 80 -255 114
rect -129 80 -113 114
rect -79 80 -63 114
rect 63 80 79 114
rect 113 80 129 114
rect 255 80 271 114
rect 305 80 321 114
rect -449 30 -415 46
rect -449 -46 -415 -30
rect -353 30 -319 46
rect -353 -46 -319 -30
rect -257 30 -223 46
rect -257 -46 -223 -30
rect -161 30 -127 46
rect -161 -46 -127 -30
rect -65 30 -31 46
rect -65 -46 -31 -30
rect 31 30 65 46
rect 31 -46 65 -30
rect 127 30 161 46
rect 127 -46 161 -30
rect 223 30 257 46
rect 223 -46 257 -30
rect 319 30 353 46
rect 319 -46 353 -30
rect 415 30 449 46
rect 415 -46 449 -30
rect -417 -114 -401 -80
rect -367 -114 -351 -80
rect -225 -114 -209 -80
rect -175 -114 -159 -80
rect -33 -114 -17 -80
rect 17 -114 33 -80
rect 159 -114 175 -80
rect 209 -114 225 -80
rect 351 -114 367 -80
rect 401 -114 417 -80
<< viali >>
rect -449 -30 -415 30
rect -353 -30 -319 30
rect -257 -30 -223 30
rect -161 -30 -127 30
rect -65 -30 -31 30
rect 31 -30 65 30
rect 127 -30 161 30
rect 223 -30 257 30
rect 319 -30 353 30
rect 415 -30 449 30
<< metal1 >>
rect -455 30 -409 42
rect -455 -30 -449 30
rect -415 -30 -409 30
rect -455 -42 -409 -30
rect -359 30 -313 42
rect -359 -30 -353 30
rect -319 -30 -313 30
rect -359 -42 -313 -30
rect -263 30 -217 42
rect -263 -30 -257 30
rect -223 -30 -217 30
rect -263 -42 -217 -30
rect -167 30 -121 42
rect -167 -30 -161 30
rect -127 -30 -121 30
rect -167 -42 -121 -30
rect -71 30 -25 42
rect -71 -30 -65 30
rect -31 -30 -25 30
rect -71 -42 -25 -30
rect 25 30 71 42
rect 25 -30 31 30
rect 65 -30 71 30
rect 25 -42 71 -30
rect 121 30 167 42
rect 121 -30 127 30
rect 161 -30 167 30
rect 121 -42 167 -30
rect 217 30 263 42
rect 217 -30 223 30
rect 257 -30 263 30
rect 217 -42 263 -30
rect 313 30 359 42
rect 313 -30 319 30
rect 353 -30 359 30
rect 313 -42 359 -30
rect 409 30 455 42
rect 409 -30 415 30
rect 449 -30 455 30
rect 409 -42 455 -30
<< properties >>
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 0.420 l 0.150 m 1 nf 9 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 0 botc 0 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 0 viasrc 100 viadrn 100 viagate 0 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
