magic
tech sky130A
magscale 1 2
timestamp 1699075837
<< error_p >>
rect 57529 57744 57537 57746
rect 57557 57744 57565 57746
rect 20103 57738 20111 57740
rect 20131 57738 20139 57740
rect 71927 57734 71935 57736
rect 71955 57734 71963 57736
rect 20095 55646 20103 55648
rect 20123 55646 20131 55648
rect 71919 55642 71927 55644
rect 71947 55642 71955 55644
rect 57499 55638 57507 55640
rect 57527 55638 57535 55640
rect 20071 53552 20079 53554
rect 20099 53552 20107 53554
rect 71895 53548 71903 53550
rect 71923 53548 71931 53550
rect 57503 53544 57511 53546
rect 57531 53544 57539 53546
<< nwell >>
rect -8858 20399 -8340 20965
<< metal1 >>
rect 103730 60470 103888 60520
rect 103730 59912 103764 60470
rect 103852 59912 103888 60470
rect 103730 59911 103888 59912
rect 103730 59877 104063 59911
rect 103730 59780 103888 59877
rect -3290 58692 -3124 58760
rect -3290 57994 -3238 58692
rect -3154 57994 -3124 58692
rect -3610 28804 -3444 28855
rect -3634 26074 -3468 26308
rect -3634 25204 -3596 26074
rect -3502 25204 -3468 26074
rect -14374 15726 -14278 15834
rect -3634 -21452 -3468 25204
rect -3290 12352 -3124 57994
rect -2970 56598 -2822 56688
rect -2970 55900 -2936 56598
rect -2852 55900 -2822 56598
rect -2970 24162 -2822 55900
rect -2330 54500 -2164 54543
rect -2330 53802 -2294 54500
rect -2210 53802 -2164 54500
rect -2970 14472 -2804 24162
rect -2970 13612 -2946 14472
rect -2852 13612 -2804 14472
rect -2970 13483 -2804 13612
rect -2650 24058 -2484 24162
rect -2650 23188 -2606 24058
rect -2512 23188 -2484 24058
rect -3290 11492 -3238 12352
rect -3144 11492 -3124 12352
rect -3290 11482 -3124 11492
rect -2650 -19328 -2484 23188
rect -2330 16540 -2164 53802
rect -1690 52400 -1524 52474
rect -1690 51702 -1638 52400
rect -1554 51702 -1524 52400
rect -2330 15680 -2284 16540
rect -2190 15680 -2164 16540
rect -2330 15647 -2164 15680
rect -2010 21994 -1844 22016
rect -2010 21124 -1976 21994
rect -1882 21124 -1844 21994
rect -2010 -17302 -1844 21124
rect -1690 18604 -1524 51702
rect -1050 50300 -884 50353
rect -1050 49602 -1002 50300
rect -918 49602 -884 50300
rect -1050 20688 -884 49602
rect -730 48222 -564 48247
rect -730 47524 -696 48222
rect -612 47524 -564 48222
rect -730 22740 -564 47524
rect -410 46134 -244 46178
rect -410 45436 -362 46134
rect -278 45436 -244 46134
rect -410 24828 -244 45436
rect -50 44034 116 44096
rect -50 43336 2 44034
rect 86 43336 116 44034
rect -50 26906 116 43336
rect 93340 31196 93476 31208
rect 93340 31164 94234 31196
rect 93340 31024 93380 31164
rect 94184 31024 94234 31164
rect 93340 31002 94234 31024
rect 93340 29082 93476 31002
rect 93290 29018 93562 29082
rect 93290 28230 93336 29018
rect 93518 28934 93562 29018
rect 93518 28230 93566 28934
rect 93290 28180 93566 28230
rect 46468 28070 46998 28113
rect 46468 27977 46830 28070
rect 46790 27288 46830 27977
rect 46956 27288 46998 28070
rect 93294 28032 93566 28180
rect 93338 28011 93474 28032
rect 46790 27256 46998 27288
rect 103750 27272 103882 59780
rect 46862 27254 46998 27256
rect -50 26140 -8 26906
rect 86 26140 116 26906
rect -50 26070 116 26140
rect -410 24062 -372 24828
rect -278 24062 -244 24828
rect -410 23982 -244 24062
rect -730 21974 -684 22740
rect -590 21974 -564 22740
rect -730 21933 -564 21974
rect -1050 19922 -1018 20688
rect -924 19922 -884 20688
rect -1690 17744 -1658 18604
rect -1564 17744 -1524 18604
rect -1690 17731 -1524 17744
rect -1370 19832 -1204 19882
rect -1370 18962 -1330 19832
rect -1236 18962 -1204 19832
rect -1050 19817 -884 19922
rect -1370 -15204 -1204 18962
rect -1050 17790 -884 17808
rect -1050 16920 -1018 17790
rect -924 16920 -884 17790
rect -1050 -13132 -884 16920
rect -730 15682 -564 15704
rect -730 14812 -696 15682
rect -602 14812 -564 15682
rect -730 -11094 -564 14812
rect -410 13618 -244 13630
rect -410 12748 -368 13618
rect -274 12748 -244 13618
rect -410 -7786 -244 12748
rect -50 11504 116 11542
rect -50 10634 -8 11504
rect 86 10634 116 11504
rect -50 -6878 116 10634
rect 23479 10298 23609 10309
rect 23352 10293 23700 10298
rect 23351 10186 23700 10293
rect 23351 9734 23400 10186
rect 22477 9676 23400 9734
rect 23662 9972 23700 10186
rect 70346 10258 70582 10362
rect 23662 9676 23710 9972
rect 70346 9758 70388 10258
rect 22477 9604 23710 9676
rect 68699 9660 70388 9758
rect 70530 9660 70582 10258
rect 68699 9628 70582 9660
rect 70346 9618 70582 9628
rect 23384 -6547 23710 9604
rect 25446 -2586 25582 -2584
rect 24478 -2646 25582 -2586
rect 24478 -2770 24544 -2646
rect 25460 -2770 25582 -2646
rect 24478 -2810 25582 -2770
rect 25446 -5811 25582 -2810
rect 71744 -5709 72066 -5690
rect 71744 -5762 72490 -5709
rect 71744 -6422 71794 -5762
rect 71994 -5845 72490 -5762
rect 71994 -6422 72066 -5845
rect 71744 -6478 72066 -6422
rect -50 -7722 -32 -6878
rect 82 -7722 116 -6878
rect -50 -7786 116 -7722
rect -410 -8918 -248 -7786
rect -410 -9762 -374 -8918
rect -260 -9208 -248 -8918
rect -260 -9762 -244 -9208
rect -410 -9908 -244 -9762
rect -730 -11938 -700 -11094
rect -586 -11938 -564 -11094
rect -730 -11960 -564 -11938
rect -1050 -13976 -1024 -13132
rect -910 -13976 -884 -13132
rect -1050 -14012 -884 -13976
rect -1370 -16048 -1334 -15204
rect -1220 -16048 -1204 -15204
rect -1370 -16092 -1204 -16048
rect -2010 -18146 -1980 -17302
rect -1866 -18146 -1844 -17302
rect -2010 -18224 -1844 -18146
rect -2650 -20172 -2632 -19328
rect -2518 -20172 -2484 -19328
rect -2650 -20388 -2484 -20172
rect -3634 -22296 -3614 -21452
rect -3500 -22296 -3468 -21452
rect -3634 -22438 -3468 -22296
rect 48266 -23530 48472 -23490
rect 95273 -23524 95403 -23521
rect 48266 -24164 48302 -23530
rect 48432 -24064 48472 -23530
rect 95270 -23574 95432 -23524
rect 48432 -24164 50627 -24064
rect 48266 -24192 50627 -24164
rect 48307 -24194 50627 -24192
rect 95270 -24204 95286 -23574
rect 95412 -24088 95432 -23574
rect 95412 -24204 97531 -24088
rect 95270 -24218 97531 -24204
rect 95270 -24234 95432 -24218
<< via1 >>
rect 103764 59912 103852 60470
rect -3238 57994 -3154 58692
rect -3596 25204 -3502 26074
rect -2936 55900 -2852 56598
rect -2294 53802 -2210 54500
rect -2946 13612 -2852 14472
rect -2606 23188 -2512 24058
rect -3238 11492 -3144 12352
rect -1638 51702 -1554 52400
rect -2284 15680 -2190 16540
rect -1976 21124 -1882 21994
rect -1002 49602 -918 50300
rect -696 47524 -612 48222
rect -362 45436 -278 46134
rect 2 43336 86 44034
rect 93380 31024 94184 31164
rect 93336 28230 93518 29018
rect 46830 27288 46956 28070
rect -8 26140 86 26906
rect -372 24062 -278 24828
rect -684 21974 -590 22740
rect -1018 19922 -924 20688
rect -1658 17744 -1564 18604
rect -1330 18962 -1236 19832
rect -1018 16920 -924 17790
rect -696 14812 -602 15682
rect -368 12748 -274 13618
rect -8 10634 86 11504
rect 23400 9676 23662 10186
rect 70388 9660 70530 10258
rect 24544 -2770 25460 -2646
rect 71794 -6422 71994 -5762
rect -32 -7722 82 -6878
rect -374 -9762 -260 -8918
rect -700 -11938 -586 -11094
rect -1024 -13976 -910 -13132
rect -1334 -16048 -1220 -15204
rect -1980 -18146 -1866 -17302
rect -2632 -20172 -2518 -19328
rect -3614 -22296 -3500 -21452
rect 48302 -24164 48432 -23530
rect 95286 -24204 95412 -23574
<< metal2 >>
rect 103518 60520 103880 60524
rect 103518 60470 103886 60520
rect 103518 60440 103764 60470
rect 103730 59912 103764 60440
rect 103852 59966 103886 60470
rect 103852 59912 104072 59966
rect 103730 59882 104072 59912
rect 103730 59878 103886 59882
rect -3278 58738 -3110 58754
rect -3299 58692 2097 58738
rect -3278 57994 -3238 58692
rect -3154 57994 -3110 58692
rect -3278 57922 -3110 57994
rect -2976 56632 -2808 56664
rect -2976 56598 2023 56632
rect -2976 55900 -2936 56598
rect -2852 56586 2023 56598
rect -2852 55900 -2808 56586
rect -2976 55832 -2808 55900
rect -2342 54538 -2174 54550
rect -3201 54500 3038 54538
rect -3201 54492 -2294 54500
rect -2342 53802 -2294 54492
rect -2210 54492 3038 54500
rect -2210 53802 -2174 54492
rect -2342 53718 -2174 53802
rect -1670 52444 -1502 52482
rect -1679 52400 2061 52444
rect -1679 52398 -1638 52400
rect -1670 51702 -1638 52398
rect -1554 52398 2061 52400
rect -1554 51702 -1502 52398
rect -1670 51650 -1502 51702
rect -1060 50350 -892 50368
rect -1060 50304 2087 50350
rect -1060 50300 -892 50304
rect -1060 49602 -1002 50300
rect -918 49602 -892 50300
rect -1060 49536 -892 49602
rect -732 48256 -564 48278
rect -733 48222 2071 48256
rect -733 48210 -696 48222
rect -732 47524 -696 48210
rect -612 48210 2071 48222
rect -612 47524 -564 48210
rect -732 47446 -564 47524
rect -408 46162 -240 46184
rect -408 46134 2111 46162
rect -408 45436 -362 46134
rect -278 46116 2111 46134
rect -278 45436 -240 46116
rect -408 45352 -240 45436
rect -50 44066 118 44096
rect -53 44034 2105 44066
rect -53 44020 2 44034
rect -50 43336 2 44020
rect 86 44020 2105 44034
rect 86 43336 118 44020
rect -50 43264 118 43336
rect 127298 42248 130768 42332
rect 93456 31196 119986 31198
rect 93340 31164 119986 31196
rect 93340 31024 93380 31164
rect 94184 31134 119986 31164
rect 94184 31024 94234 31134
rect 93340 31002 94234 31024
rect 93340 29082 93476 31002
rect 93290 29018 93562 29082
rect 93290 28230 93336 29018
rect 93518 28230 93562 29018
rect 93290 28180 93562 28230
rect 46790 28070 46994 28112
rect 46790 27288 46830 28070
rect 46956 27397 46994 28070
rect 119922 27423 119986 31134
rect 130684 27423 130768 42248
rect 46956 27333 48948 27397
rect 116760 27359 130792 27423
rect 46956 27288 46994 27333
rect 46790 27256 46994 27288
rect -44 26906 122 27000
rect -44 26140 -8 26906
rect 86 26140 122 26906
rect -44 26130 122 26140
rect -6742 26082 1758 26130
rect -7646 22438 -7188 22450
rect -6742 22438 -6694 26082
rect -3634 26074 -3458 26082
rect -44 26074 122 26082
rect -3634 25204 -3596 26074
rect -3502 25204 -3458 26074
rect -3634 25146 -3458 25204
rect -404 24828 -238 24932
rect -2644 24058 -2468 24112
rect -2644 24044 -2606 24058
rect -7646 22416 -6694 22438
rect -8014 22414 -6694 22416
rect -8014 22354 -7960 22414
rect -7260 22390 -6694 22414
rect -6220 23996 -2606 24044
rect -7260 22354 -7188 22390
rect -8014 22320 -7188 22354
rect -8018 21314 -7192 21364
rect -8018 21254 -7970 21314
rect -7270 21306 -7192 21314
rect -6220 21306 -6172 23996
rect -2644 23188 -2606 23996
rect -2512 24044 -2468 24058
rect -404 24062 -372 24828
rect -278 24062 -238 24828
rect -404 24044 -238 24062
rect -2512 23996 1760 24044
rect -2512 23188 -2468 23996
rect -2644 23150 -2468 23188
rect -726 22740 -560 22848
rect -2008 21994 -1832 22040
rect -2008 21950 -1976 21994
rect -7270 21258 -6172 21306
rect -5766 21902 -1976 21950
rect -7270 21254 -7192 21258
rect -8018 21234 -7192 21254
rect -7994 20230 -7168 20274
rect -7994 20170 -7954 20230
rect -7254 20208 -7168 20230
rect -5766 20208 -5718 21902
rect -2008 21124 -1976 21902
rect -1882 21950 -1832 21994
rect -726 21974 -684 22740
rect -590 21974 -560 22740
rect -726 21950 -560 21974
rect -1882 21902 1726 21950
rect -1882 21124 -1832 21902
rect -2008 21078 -1832 21124
rect -7254 20170 -5718 20208
rect -7994 20160 -5718 20170
rect -7994 20144 -7168 20160
rect -5766 20150 -5718 20160
rect -1044 20688 -878 20764
rect -1044 19922 -1018 20688
rect -924 19922 -878 20688
rect -1382 19860 -1206 19868
rect -1044 19860 -878 19922
rect -7096 19832 1786 19860
rect -7096 19812 -1330 19832
rect -8018 19144 -7192 19184
rect -8018 19084 -7970 19144
rect -7270 19134 -7192 19144
rect -7096 19134 -7048 19812
rect -7270 19086 -7048 19134
rect -7270 19084 -7192 19086
rect -8018 19054 -7192 19084
rect -1382 18962 -1330 19812
rect -1236 19812 1786 19832
rect -1236 18962 -1206 19812
rect -1382 18906 -1206 18962
rect -1700 18604 -1534 18648
rect -7998 18090 -4354 18124
rect -8028 18076 -4354 18090
rect -8028 18064 -7202 18076
rect -8028 18004 -7954 18064
rect -7254 18004 -7202 18064
rect -8028 17960 -7202 18004
rect -4402 17762 -4354 18076
rect -1700 17762 -1658 18604
rect -4402 17744 -1658 17762
rect -1564 17762 -1534 18604
rect -1060 17790 -884 17810
rect -1060 17762 -1018 17790
rect -1564 17744 -1018 17762
rect -4402 17714 -1018 17744
rect -8004 16974 -7178 17004
rect -8004 16914 -7954 16974
rect -7254 16972 -7178 16974
rect -7254 16924 -4732 16972
rect -7254 16914 -7178 16924
rect -8004 16874 -7178 16914
rect -8012 15892 -5630 15940
rect -8008 15874 -7182 15892
rect -8008 15814 -7960 15874
rect -7260 15814 -7182 15874
rect -8008 15788 -7182 15814
rect -8018 14810 -7086 14818
rect -8018 14798 -6628 14810
rect -8018 14724 -7964 14798
rect -7270 14762 -6628 14798
rect -7270 14724 -7086 14762
rect -8018 14704 -7086 14724
rect -6676 11500 -6628 14762
rect -5678 13586 -5630 15892
rect -4780 15680 -4732 16924
rect -1060 16920 -1018 17714
rect -924 17762 -884 17790
rect -924 17714 1846 17762
rect -924 16920 -884 17714
rect -1060 16848 -884 16920
rect -2320 16540 -2154 16566
rect -2320 15680 -2284 16540
rect -2190 15680 -2154 16540
rect -742 15682 -566 15726
rect -742 15680 -696 15682
rect -4780 15632 -696 15680
rect -742 14812 -696 15632
rect -602 15680 -566 15682
rect -602 15632 1832 15680
rect -602 14812 -566 15632
rect -742 14764 -566 14812
rect -2972 13612 -2946 14472
rect -2852 13612 -2806 14472
rect -2972 13586 -2806 13612
rect -398 13618 -222 13658
rect -398 13586 -368 13618
rect -5678 13538 -368 13586
rect -398 12748 -368 13538
rect -274 13586 -222 13618
rect -274 13538 1782 13586
rect -274 12748 -222 13538
rect -398 12696 -222 12748
rect -3278 12352 -3112 12398
rect -3278 11500 -3238 12352
rect -6676 11492 -3238 11500
rect -3144 11500 -3112 12352
rect -54 11504 122 11544
rect -54 11500 -8 11504
rect -3144 11492 -8 11500
rect -6676 11452 -8 11492
rect -54 10634 -8 11452
rect 86 11500 122 11504
rect 86 11452 1844 11500
rect 86 10634 122 11452
rect -54 10582 122 10634
rect 70346 10329 70582 10362
rect 23352 10295 23700 10298
rect 23352 10186 25455 10295
rect 3494 -2580 3734 9747
rect 23352 9676 23400 10186
rect 23662 10181 25455 10186
rect 70346 10258 72813 10329
rect 23662 9676 23700 10181
rect 23352 9618 23700 9676
rect 70346 9660 70388 10258
rect 70530 10215 72813 10258
rect 70530 9660 70582 10215
rect 70346 9618 70582 9660
rect 3494 -2646 25606 -2580
rect 3494 -2770 24544 -2646
rect 25460 -2770 25606 -2646
rect 3494 -2820 25606 -2770
rect 3494 -6524 3734 -2820
rect 71744 -5762 72066 -5690
rect 71744 -6422 71794 -5762
rect 71994 -6422 72066 -5762
rect 71744 -6425 72066 -6422
rect 70558 -6478 72066 -6425
rect 70558 -6489 72010 -6478
rect -64 -6878 132 -6808
rect -64 -7722 -32 -6878
rect 82 -7681 132 -6878
rect 82 -7722 3062 -7681
rect -64 -7729 3062 -7722
rect -64 -7758 132 -7729
rect -410 -8918 -214 -8880
rect -410 -9762 -374 -8918
rect -260 -9762 -214 -8918
rect -410 -9767 -214 -9762
rect -410 -9815 3046 -9767
rect -410 -9830 -214 -9815
rect -750 -11094 -554 -11020
rect -750 -11938 -700 -11094
rect -586 -11861 -554 -11094
rect -586 -11909 3030 -11861
rect -586 -11938 -554 -11909
rect -750 -11970 -554 -11938
rect -1066 -13132 -870 -13066
rect -1066 -13976 -1024 -13132
rect -910 -13951 -870 -13132
rect -910 -13976 3128 -13951
rect -1066 -13999 3128 -13976
rect -1066 -14016 -870 -13999
rect -1382 -15204 -1186 -15150
rect -1382 -16048 -1334 -15204
rect -1220 -16048 -1186 -15204
rect -1382 -16049 -1186 -16048
rect -1382 -16092 3122 -16049
rect -1382 -16100 -1186 -16092
rect -876 -16097 3122 -16092
rect -2018 -17302 -1822 -17252
rect -2018 -18146 -1980 -17302
rect -1866 -18131 -1822 -17302
rect -1866 -18146 3106 -18131
rect -2018 -18179 3106 -18146
rect -2018 -18202 -1822 -18179
rect -2668 -19328 -2472 -19294
rect -2668 -20172 -2632 -19328
rect -2518 -20172 -2472 -19328
rect -2668 -20225 -2472 -20172
rect -2668 -20244 3134 -20225
rect -2636 -20273 3134 -20244
rect -3656 -21452 -3460 -21366
rect -3656 -22296 -3614 -21452
rect -3500 -22296 -3460 -21452
rect -3656 -22311 -3460 -22296
rect -3656 -22316 3118 -22311
rect -3630 -22359 3118 -22316
rect 48266 -23493 48472 -23490
rect 45511 -23530 48473 -23493
rect 95270 -23527 95432 -23524
rect 45511 -23607 48302 -23530
rect 48266 -24164 48302 -23607
rect 48432 -23607 48473 -23530
rect 92875 -23574 95432 -23527
rect 48432 -24164 48472 -23607
rect 92875 -23641 95286 -23574
rect 48266 -24192 48472 -24164
rect 95270 -24204 95286 -23641
rect 95412 -24204 95432 -23574
rect 95270 -24234 95432 -24204
<< via2 >>
rect -7960 22354 -7260 22414
rect -7970 21254 -7270 21314
rect -7954 20170 -7254 20230
rect -7970 19084 -7270 19144
rect -7954 18004 -7254 18064
rect -7954 16914 -7254 16974
rect -7960 15814 -7260 15874
rect -7964 14724 -7270 14798
<< metal3 >>
rect -6135 33318 -5077 33329
rect -6139 32940 6171 33318
rect -6135 309 -5077 32940
rect -6156 -83 3438 309
rect -6135 -33083 -5077 -83
rect -6135 -34141 6745 -33083
<< metal4 >>
rect 117713 26377 118267 34013
rect 378 24503 421 25057
rect -14447 21912 -14127 22416
rect -12745 15738 -12425 16092
rect -10383 13176 -10063 16138
rect -9341 14657 -9021 17040
rect -9341 14122 449 14657
rect -8424 14103 449 14122
rect -10383 13034 -8348 13176
rect -10383 12652 -10274 13034
rect -8458 12652 -8348 13034
rect -10383 12628 -8348 12652
rect -10338 12604 -8348 12628
rect 117253 -7029 117951 1024
<< via4 >>
rect -10274 12652 -8458 13034
<< metal5 >>
rect 378 25129 556 25701
rect 118220 24658 118792 33044
rect -14124 21998 -13804 22416
rect -10353 13034 559 13151
rect -10353 12652 -10274 13034
rect -8458 12652 559 13034
rect -10353 12597 559 12652
rect 118220 -6080 118792 262
use cp1_buffer_5stage  cp1_buffer_5stage_0
timestamp 1699075837
transform 1 0 58 0 1 32336
box -1331 -130 130524 30508
use cp2_buffer_5stage  cp2_buffer_5stage_0
timestamp 1699074715
transform -1 0 93962 0 1 -1060
box -25261 108 95113 31581
use cp2_buffer_5stage  cp2_buffer_5stage_1
timestamp 1699074715
transform 1 0 24944 0 1 -34882
box -25261 108 95113 31581
use scanchain  scanchain_0
timestamp 1698771642
transform 1 0 -16242 0 1 13610
box 158 1096 9026 9920
<< end >>
