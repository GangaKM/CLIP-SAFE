magic
tech sky130A
magscale 1 2
timestamp 1698753667
<< nwell >>
rect 768 15858 974 15860
rect 768 15530 976 15858
rect 780 15132 976 15530
rect 24064 7868 24318 8204
<< psubdiff >>
rect 18057 18772 21688 18848
rect 3340 18612 7634 18650
rect 3340 18152 3472 18612
rect 7492 18152 7634 18612
rect 18057 18340 18164 18772
rect 21510 18340 21688 18772
rect 18057 18271 21688 18340
rect 3340 18086 7634 18152
<< nsubdiff >>
rect 12396 17402 12508 17434
rect 12396 17294 12430 17402
rect 12484 17294 12508 17402
rect 12396 17274 12508 17294
rect 840 15788 934 15820
rect 840 15546 860 15788
rect 916 15546 934 15788
rect 840 15520 934 15546
rect 24100 8124 24242 8162
rect 24100 7934 24128 8124
rect 24206 7934 24242 8124
rect 24100 7904 24242 7934
<< psubdiffcont >>
rect 3472 18152 7492 18612
rect 18164 18340 21510 18772
<< nsubdiffcont >>
rect 12430 17294 12484 17402
rect 860 15546 916 15788
rect 24128 7934 24206 8124
<< poly >>
rect 24310 16424 24438 16600
rect 24310 16394 24468 16424
rect 24310 16232 24438 16394
rect 24310 16202 24490 16232
rect 24310 16040 24438 16202
rect 24310 16010 24488 16040
rect 24310 15848 24438 16010
rect 402 15666 584 15824
rect 402 15636 628 15666
rect 402 15474 584 15636
rect 24310 15818 24488 15848
rect 24310 15656 24438 15818
rect 24310 15626 24486 15656
rect 402 15444 634 15474
rect 24310 15464 24438 15626
rect 402 15282 584 15444
rect 24310 15434 24476 15464
rect 402 15252 632 15282
rect 24310 15272 24438 15434
rect 402 15090 584 15252
rect 24310 15242 24480 15272
rect 402 15060 630 15090
rect 24310 15080 24438 15242
rect 402 14898 584 15060
rect 24310 15050 24464 15080
rect 402 14868 626 14898
rect 24310 14888 24438 15050
rect 402 14706 584 14868
rect 24310 14858 24466 14888
rect 402 14676 632 14706
rect 24310 14696 24438 14858
rect 402 14514 584 14676
rect 24310 14666 24476 14696
rect 402 14484 630 14514
rect 24310 14504 24438 14666
rect 402 14322 584 14484
rect 24310 14474 24472 14504
rect 402 14292 632 14322
rect 24310 14312 24438 14474
rect 402 14130 584 14292
rect 24310 14282 24470 14312
rect 402 14100 632 14130
rect 24310 14120 24438 14282
rect 402 13938 584 14100
rect 24310 14090 24478 14120
rect 402 13908 632 13938
rect 24310 13928 24438 14090
rect 402 13746 584 13908
rect 24310 13898 24478 13928
rect 402 13716 642 13746
rect 24310 13736 24438 13898
rect 402 13554 584 13716
rect 24310 13706 24476 13736
rect 402 13524 638 13554
rect 24310 13544 24438 13706
rect 402 13362 584 13524
rect 24310 13514 24466 13544
rect 402 13332 632 13362
rect 24310 13352 24438 13514
rect 402 13170 584 13332
rect 24310 13322 24480 13352
rect 402 13140 630 13170
rect 24310 13160 24438 13322
rect 402 12978 584 13140
rect 24310 13130 24474 13160
rect 402 12948 632 12978
rect 24310 12968 24438 13130
rect 402 12786 584 12948
rect 24310 12938 24474 12968
rect 402 12756 640 12786
rect 24310 12776 24438 12938
rect 402 12594 584 12756
rect 24310 12746 24470 12776
rect 402 12564 628 12594
rect 24310 12584 24438 12746
rect 402 12402 584 12564
rect 24310 12554 24478 12584
rect 402 12372 630 12402
rect 24310 12392 24438 12554
rect 402 12210 584 12372
rect 24310 12362 24472 12392
rect 402 12180 636 12210
rect 24310 12200 24438 12362
rect 402 12018 584 12180
rect 24310 12170 24478 12200
rect 402 11988 632 12018
rect 24310 12008 24438 12170
rect 402 11826 584 11988
rect 24310 11978 24470 12008
rect 402 11796 628 11826
rect 24310 11816 24438 11978
rect 402 11634 584 11796
rect 24310 11786 24472 11816
rect 402 11604 630 11634
rect 24310 11624 24438 11786
rect 402 11442 584 11604
rect 24310 11594 24470 11624
rect 402 11412 626 11442
rect 24310 11432 24438 11594
rect 402 11250 584 11412
rect 24310 11402 24478 11432
rect 402 11220 632 11250
rect 24310 11240 24438 11402
rect 402 11058 584 11220
rect 24310 11210 24474 11240
rect 402 11028 642 11058
rect 24310 11048 24438 11210
rect 402 10866 584 11028
rect 24310 11018 24476 11048
rect 402 10836 630 10866
rect 24310 10856 24438 11018
rect 402 10674 584 10836
rect 24310 10826 24476 10856
rect 402 10644 638 10674
rect 24310 10664 24438 10826
rect 402 10482 584 10644
rect 24310 10634 24480 10664
rect 402 10452 640 10482
rect 24310 10472 24438 10634
rect 402 10290 584 10452
rect 24310 10442 24474 10472
rect 402 10260 634 10290
rect 24310 10280 24438 10442
rect 402 10098 584 10260
rect 24310 10250 24476 10280
rect 402 10068 626 10098
rect 24310 10088 24438 10250
rect 402 9906 584 10068
rect 24310 10058 24476 10088
rect 402 9876 630 9906
rect 24310 9896 24438 10058
rect 402 9714 584 9876
rect 24310 9866 24484 9896
rect 402 9684 632 9714
rect 24310 9704 24438 9866
rect 402 9522 584 9684
rect 24310 9674 24460 9704
rect 402 9492 634 9522
rect 24310 9512 24438 9674
rect 402 9330 584 9492
rect 24310 9482 24476 9512
rect 402 9300 634 9330
rect 24310 9320 24438 9482
rect 402 9138 584 9300
rect 24310 9290 24468 9320
rect 402 9108 632 9138
rect 24310 9128 24438 9290
rect 402 8946 584 9108
rect 24310 9098 24466 9128
rect 402 8916 626 8946
rect 24310 8936 24438 9098
rect 402 8754 584 8916
rect 24310 8908 24478 8936
rect 24422 8906 24478 8908
rect 402 8724 626 8754
rect 402 8562 584 8724
rect 402 8532 628 8562
rect 402 8370 584 8532
rect 402 8340 634 8370
rect 402 8178 584 8340
rect 402 8148 632 8178
rect 402 8144 584 8148
rect 24500 8102 24560 8218
rect 24468 8072 24560 8102
rect 636 7918 702 7926
rect 614 7888 702 7918
rect 24500 7910 24560 8072
rect 636 7726 702 7888
rect 24472 7880 24560 7910
rect 612 7696 702 7726
rect 24500 7718 24560 7880
rect 636 7534 702 7696
rect 24476 7688 24560 7718
rect 610 7504 702 7534
rect 24500 7526 24560 7688
rect 636 7342 702 7504
rect 24468 7496 24560 7526
rect 610 7312 702 7342
rect 24500 7334 24560 7496
rect 636 7150 702 7312
rect 24470 7304 24560 7334
rect 612 7120 702 7150
rect 24500 7142 24560 7304
rect 636 6958 702 7120
rect 24472 7112 24560 7142
rect 614 6928 702 6958
rect 24500 6950 24560 7112
rect 636 6766 702 6928
rect 24472 6920 24560 6950
rect 610 6736 702 6766
rect 24500 6758 24560 6920
rect 636 6574 702 6736
rect 24470 6728 24560 6758
rect 610 6544 702 6574
rect 24500 6566 24560 6728
rect 636 6382 702 6544
rect 24472 6536 24560 6566
rect 612 6352 702 6382
rect 24500 6374 24560 6536
rect 636 6190 702 6352
rect 24476 6344 24560 6374
rect 610 6160 702 6190
rect 24500 6182 24560 6344
rect 636 5998 702 6160
rect 24476 6152 24560 6182
rect 612 5968 702 5998
rect 24500 5990 24560 6152
rect 636 5806 702 5968
rect 24476 5960 24560 5990
rect 612 5776 702 5806
rect 24500 5798 24560 5960
rect 636 5614 702 5776
rect 24470 5768 24560 5798
rect 612 5584 702 5614
rect 24500 5606 24560 5768
rect 636 5422 702 5584
rect 24470 5576 24560 5606
rect 614 5392 702 5422
rect 24500 5414 24560 5576
rect 636 5230 702 5392
rect 24476 5384 24560 5414
rect 610 5200 702 5230
rect 24500 5222 24560 5384
rect 636 5038 702 5200
rect 24470 5192 24560 5222
rect 608 5008 702 5038
rect 24500 5030 24560 5192
rect 636 4846 702 5008
rect 24472 5000 24560 5030
rect 610 4816 702 4846
rect 24500 4838 24560 5000
rect 636 4654 702 4816
rect 24472 4808 24560 4838
rect 612 4624 702 4654
rect 24500 4646 24560 4808
rect 636 4462 702 4624
rect 24468 4616 24560 4646
rect 610 4432 702 4462
rect 24500 4454 24560 4616
rect 636 4270 702 4432
rect 24474 4424 24560 4454
rect 612 4240 702 4270
rect 24500 4262 24560 4424
rect 636 4078 702 4240
rect 24472 4232 24560 4262
rect 610 4048 702 4078
rect 24500 4070 24560 4232
rect 636 3886 702 4048
rect 24470 4040 24560 4070
rect 614 3856 702 3886
rect 24500 3878 24560 4040
rect 636 3694 702 3856
rect 24472 3848 24560 3878
rect 612 3664 702 3694
rect 24500 3686 24560 3848
rect 636 3502 702 3664
rect 24472 3656 24560 3686
rect 616 3472 702 3502
rect 24500 3494 24560 3656
rect 636 3310 702 3472
rect 24474 3464 24560 3494
rect 612 3280 702 3310
rect 24500 3302 24560 3464
rect 636 3118 702 3280
rect 24470 3272 24560 3302
rect 618 3088 702 3118
rect 24500 3110 24560 3272
rect 636 2926 702 3088
rect 24472 3080 24560 3110
rect 612 2896 702 2926
rect 24500 2918 24560 3080
rect 636 2734 702 2896
rect 24476 2888 24560 2918
rect 616 2704 702 2734
rect 24500 2726 24560 2888
rect 636 2542 702 2704
rect 24472 2696 24560 2726
rect 614 2512 702 2542
rect 24500 2534 24560 2696
rect 636 2350 702 2512
rect 24474 2504 24560 2534
rect 614 2320 702 2350
rect 24500 2342 24560 2504
rect 636 2158 702 2320
rect 24466 2312 24560 2342
rect 616 2128 702 2158
rect 24500 2150 24560 2312
rect 636 1966 702 2128
rect 24472 2120 24560 2150
rect 614 1936 702 1966
rect 24500 1958 24560 2120
rect 636 1774 702 1936
rect 24474 1928 24560 1958
rect 618 1744 702 1774
rect 24500 1766 24560 1928
rect 636 1582 702 1744
rect 24476 1736 24560 1766
rect 616 1552 702 1582
rect 24500 1574 24560 1736
rect 636 1390 702 1552
rect 24472 1544 24560 1574
rect 616 1360 702 1390
rect 24500 1382 24560 1544
rect 636 1198 702 1360
rect 24468 1352 24560 1382
rect 614 1168 702 1198
rect 24500 1190 24560 1352
rect 636 1006 702 1168
rect 24474 1160 24560 1190
rect 622 976 702 1006
rect 24500 998 24560 1160
rect 636 814 702 976
rect 24466 968 24560 998
rect 614 784 702 814
rect 24500 806 24560 968
rect 636 622 702 784
rect 24478 776 24560 806
rect 618 592 702 622
rect 24500 614 24560 776
rect 636 430 702 592
rect 24472 584 24560 614
rect 24500 462 24560 584
rect 616 400 702 430
rect 636 230 702 400
<< locali >>
rect 18057 18772 21688 18848
rect 3340 18612 7634 18650
rect 3340 18152 3472 18612
rect 7492 18152 7634 18612
rect 18057 18340 18164 18772
rect 21510 18340 21688 18772
rect 18057 18271 21688 18340
rect 3340 18086 7634 18152
rect 12396 17402 12506 17436
rect 12396 17294 12430 17402
rect 12484 17294 12506 17402
rect 12396 17262 12506 17294
rect 24126 16486 24438 16600
rect 66 15702 584 15848
rect 66 8214 164 15702
rect 440 8214 584 15702
rect 840 15788 934 15820
rect 840 15546 860 15788
rect 916 15546 934 15788
rect 840 15520 934 15546
rect 24126 9030 24200 16486
rect 24330 9030 24438 16486
rect 24126 8908 24438 9030
rect 24126 8896 24372 8908
rect 66 8110 584 8214
rect 24502 8172 25032 8338
rect 24100 8124 24242 8162
rect 24100 7934 24128 8124
rect 24206 7934 24242 8124
rect 646 7804 1088 7930
rect 24100 7904 24242 7934
rect 646 328 806 7804
rect 1032 328 1088 7804
rect 24502 474 24732 8172
rect 24954 474 25032 8172
rect 24502 390 25032 474
rect 646 230 1088 328
<< viali >>
rect 3472 18152 7492 18612
rect 18164 18340 21510 18772
rect 12430 17294 12484 17402
rect 164 8214 440 15702
rect 860 15546 916 15788
rect 24200 9030 24330 16486
rect 24128 7934 24206 8124
rect 806 328 1032 7804
rect 24732 474 24954 8172
<< metal1 >>
rect 12684 19366 12720 19520
rect 12826 19374 12860 19517
rect 21978 19374 23760 19382
rect 944 19270 12723 19366
rect 12826 19359 23843 19374
rect 12826 19325 23887 19359
rect 944 19070 1024 19270
rect 2602 19070 12723 19270
rect 944 19036 12723 19070
rect 12832 19306 23843 19325
rect 12832 19126 22184 19306
rect 23678 19126 23843 19306
rect 12832 19060 23843 19126
rect 18057 18807 21688 18848
rect 18057 18772 24844 18807
rect 3340 18612 7634 18650
rect 3340 18493 3472 18612
rect 122 18152 3472 18493
rect 7492 18152 7634 18612
rect 18057 18340 18164 18772
rect 21510 18453 24844 18772
rect 21510 18340 21688 18453
rect 11282 18322 11684 18340
rect 11282 18282 11358 18322
rect 10696 18188 11358 18282
rect 11654 18282 11684 18322
rect 13378 18298 13984 18324
rect 13378 18288 13410 18298
rect 11654 18188 12138 18282
rect 12846 18214 13410 18288
rect 13932 18288 13984 18298
rect 13932 18214 14814 18288
rect 18057 18271 21688 18340
rect 12846 18196 14814 18214
rect 11282 18160 11684 18188
rect 13378 18182 13984 18196
rect 122 18103 7634 18152
rect 122 15702 512 18103
rect 3340 18086 7634 18103
rect 12370 18132 12534 18148
rect 12370 17290 12400 18132
rect 12502 17290 12534 18132
rect 14430 17600 14534 17698
rect 14430 17508 14720 17600
rect 12370 17240 12534 17290
rect 122 8214 164 15702
rect 440 8214 512 15702
rect 122 8170 512 8214
rect 630 16389 2043 16823
rect 24126 16486 24372 16600
rect 24126 16466 24200 16486
rect 23146 16400 24200 16466
rect 630 15788 1064 16389
rect 630 15546 860 15788
rect 916 15546 1064 15788
rect 122 8168 548 8170
rect 226 7998 548 8168
rect 630 8026 1064 15546
rect 24126 14554 24200 16400
rect 22540 14414 24200 14554
rect 24126 9030 24200 14414
rect 24330 9030 24372 16486
rect 24126 8896 24372 9030
rect 24490 15858 24844 18453
rect 24490 8810 24954 15858
rect 24732 8336 24954 8810
rect 23978 8190 24458 8232
rect 22662 8124 24458 8190
rect 22662 8086 24128 8124
rect 226 186 594 7998
rect 700 7804 1142 7936
rect 700 328 806 7804
rect 1032 6184 1142 7804
rect 23978 7934 24128 8086
rect 24206 7934 24458 8124
rect 1032 5984 2306 6184
rect 1032 2014 1142 5984
rect 1032 1788 2412 2014
rect 1032 328 1142 1788
rect 700 236 1142 328
rect 12659 300 13345 366
rect 23978 330 24458 7934
rect 24630 8172 25012 8336
rect 24630 474 24732 8172
rect 24954 474 25012 8172
rect 24630 392 25012 474
rect 10333 174 12352 252
rect 1980 108 7148 150
rect 2596 68 7148 108
rect 2596 -90 9480 68
rect 2596 -238 2720 -90
rect 3848 -238 9480 -90
rect 2596 -298 9480 -238
rect 4348 -344 4900 -326
rect 4348 -441 4368 -344
rect 4341 -494 4368 -441
rect 4880 -441 4900 -344
rect 10333 -441 10411 174
rect 4880 -494 10411 -441
rect 4341 -519 10411 -494
rect 12464 -472 12478 -410
rect 12538 -472 12550 -410
rect 12464 -576 12550 -472
rect 13279 -453 13345 300
rect 20752 154 22362 180
rect 22738 154 23106 180
rect 15520 30 17650 68
rect 20752 30 23106 154
rect 15520 -88 23106 30
rect 15520 -216 21968 -88
rect 22960 -216 23106 -88
rect 15520 -268 23106 -216
rect 20066 -442 20476 -408
rect 20066 -453 20098 -442
rect 13279 -504 20098 -453
rect 20442 -504 20476 -442
rect 13279 -519 20476 -504
rect 20066 -530 20476 -519
rect 936 -701 1482 -688
rect 8366 -701 8664 -698
rect 936 -735 10736 -701
rect 23632 -706 24074 -694
rect 936 -788 1482 -735
rect 936 -1984 1006 -788
rect 1406 -1984 1482 -788
rect 8366 -744 8664 -735
rect 14458 -742 24074 -706
rect 8366 -1102 8398 -744
rect 8632 -1102 8664 -744
rect 8366 -1446 8664 -1102
rect 16224 -750 16610 -742
rect 16224 -1082 16268 -750
rect 16572 -1082 16610 -750
rect 16224 -1464 16610 -1082
rect 23632 -752 24074 -742
rect 23632 -1826 23696 -752
rect 23998 -1826 24074 -752
rect 23632 -1902 24074 -1826
rect 936 -2064 1482 -1984
<< via1 >>
rect 1024 19070 2602 19270
rect 22184 19126 23678 19306
rect 3472 18152 7492 18612
rect 18164 18340 21510 18772
rect 11358 18188 11654 18322
rect 13410 18214 13932 18298
rect 12400 17402 12502 18132
rect 12400 17294 12430 17402
rect 12430 17294 12484 17402
rect 12484 17294 12502 17402
rect 12400 17290 12502 17294
rect 2720 -238 3848 -90
rect 4368 -494 4880 -344
rect 12478 -472 12538 -410
rect 21968 -216 22960 -88
rect 20098 -504 20442 -442
rect 1006 -1984 1406 -788
rect 8398 -1102 8632 -744
rect 16268 -1082 16572 -750
rect 23696 -1826 23998 -752
<< metal2 >>
rect 942 19270 2738 19362
rect 942 19070 1024 19270
rect 2602 19070 2738 19270
rect 942 19006 2738 19070
rect 21978 19306 23760 19382
rect 21978 19126 22184 19306
rect 23678 19126 23760 19306
rect 21978 19062 23760 19126
rect 18057 18772 21688 18848
rect 3340 18612 7634 18650
rect 3340 18152 3472 18612
rect 7492 18152 7634 18612
rect 18057 18340 18164 18772
rect 21510 18340 21688 18772
rect 11282 18322 11684 18340
rect 11282 18188 11358 18322
rect 11654 18188 11684 18322
rect 11282 18160 11684 18188
rect 13378 18298 13984 18324
rect 13378 18214 13410 18298
rect 13932 18214 13984 18298
rect 18057 18271 21688 18340
rect 13378 18182 13984 18214
rect 3340 18086 7634 18152
rect 12370 18132 12540 18174
rect 12370 17368 12400 18132
rect 12368 17290 12400 17368
rect 12502 17290 12540 18132
rect 12368 17240 12540 17290
rect 12368 17147 12534 17240
rect -313 16981 25321 17147
rect 11684 15874 13378 15926
rect 11736 13780 13362 13832
rect 11744 11696 13374 11748
rect 11720 9610 13416 9662
rect 11746 7524 13420 7576
rect 11726 5438 13352 5490
rect 11754 3354 13390 3406
rect 11662 1220 13430 1272
rect 2624 -90 3956 -46
rect 2624 -238 2720 -90
rect 3848 -238 3956 -90
rect 2624 -288 3956 -238
rect 21882 -88 23078 -40
rect 21882 -216 21968 -88
rect 22960 -216 23078 -88
rect 21882 -248 23078 -216
rect 4348 -344 4900 -326
rect 4348 -494 4368 -344
rect 4880 -494 4900 -344
rect 4348 -512 4900 -494
rect 12470 -472 12478 -410
rect 12538 -472 12550 -410
rect 12470 -534 12550 -472
rect 20066 -442 20476 -408
rect 20066 -504 20098 -442
rect 20442 -504 20476 -442
rect 20066 -530 20476 -504
rect 12466 -568 12550 -534
rect 346 -652 25164 -568
rect 936 -788 1482 -688
rect 936 -1984 1006 -788
rect 1406 -1984 1482 -788
rect 8366 -744 8664 -698
rect 8366 -1102 8398 -744
rect 8632 -1102 8664 -744
rect 8366 -1446 8664 -1102
rect 16224 -750 16610 -706
rect 16224 -1082 16268 -750
rect 16572 -1082 16610 -750
rect 16224 -1464 16610 -1082
rect 23632 -752 24074 -694
rect 23632 -1826 23696 -752
rect 23998 -1826 24074 -752
rect 23632 -1902 24074 -1826
rect 936 -2064 1482 -1984
<< via2 >>
rect 1024 19070 2602 19270
rect 22184 19126 23678 19306
rect 3472 18152 7492 18612
rect 18164 18340 21510 18772
rect 11358 18188 11654 18322
rect 13410 18214 13932 18298
rect 2720 -238 3848 -90
rect 21968 -216 22960 -88
rect 4368 -494 4880 -344
rect 20098 -504 20442 -442
rect 1006 -1984 1406 -788
rect 8398 -1102 8632 -744
rect 16268 -1082 16572 -750
rect 23696 -1826 23998 -752
<< metal3 >>
rect 944 19362 1468 19402
rect 21978 19371 23760 19382
rect 942 19270 2738 19362
rect 942 19070 1024 19270
rect 2602 19070 2738 19270
rect 942 19006 2738 19070
rect 21978 19306 24060 19371
rect 21978 19126 22184 19306
rect 23678 19126 24060 19306
rect 21978 19062 24060 19126
rect 944 17800 1468 19006
rect 18057 18772 21688 18848
rect 3340 18612 7634 18650
rect 3340 18152 3472 18612
rect 7492 18152 7634 18612
rect 18057 18340 18164 18772
rect 21510 18340 21688 18772
rect 11318 18322 11684 18340
rect 11318 18188 11358 18322
rect 11654 18188 11684 18322
rect 11318 18160 11684 18188
rect 13378 18298 13984 18324
rect 13378 18214 13410 18298
rect 13932 18214 13984 18298
rect 18057 18271 21688 18340
rect 13378 18182 13984 18214
rect 3340 18086 7634 18152
rect 23638 17970 24060 19062
rect 23502 17966 24060 17970
rect 944 17280 10212 17800
rect 944 17276 1592 17280
rect 944 1099 1464 17276
rect 12066 15806 12180 17765
rect 12714 15813 12828 17841
rect 15074 17546 24060 17966
rect 12910 15813 13417 15815
rect 11658 15805 12314 15806
rect 11658 15542 12400 15805
rect 12714 15573 13417 15813
rect 12714 15569 13244 15573
rect 11874 13734 12400 15542
rect 11364 13710 12400 13734
rect 11426 13470 12400 13710
rect 11874 11648 12400 13470
rect 11699 11402 12400 11648
rect 11874 9562 12400 11402
rect 11689 9316 12400 9562
rect 11874 7476 12400 9316
rect 11755 7230 12400 7476
rect 11874 5392 12400 7230
rect 11724 5146 12400 5392
rect 11874 3308 12400 5146
rect 11741 3062 12400 3308
rect 11874 1236 12400 3062
rect 11620 1216 12400 1236
rect 11224 1124 12400 1216
rect 944 1062 2019 1099
rect 944 1010 2033 1062
rect 11569 1058 12400 1124
rect 12718 13724 13244 15569
rect 12718 13478 13477 13724
rect 12718 11638 13244 13478
rect 12718 11392 13403 11638
rect 12718 9552 13244 11392
rect 12718 9306 13389 9552
rect 12718 7466 13244 9306
rect 12718 7220 13407 7466
rect 12718 5382 13244 7220
rect 12718 5136 13455 5382
rect 12718 1186 13244 5136
rect 13412 1186 13950 1226
rect 12718 1058 13950 1186
rect 23638 1092 24060 17546
rect 22984 1060 24060 1092
rect 944 1009 2019 1010
rect 944 -788 1464 1009
rect 2624 -90 3956 -46
rect 2624 -238 2720 -90
rect 3848 -238 3956 -90
rect 2624 -288 3956 -238
rect 4348 -344 4900 -326
rect 4348 -494 4368 -344
rect 4880 -494 4900 -344
rect 4348 -512 4900 -494
rect 944 -1984 1006 -788
rect 1406 -1984 1464 -788
rect 8368 -744 8662 -694
rect 8368 -1102 8398 -744
rect 8632 -1102 8662 -744
rect 8368 -1152 8662 -1102
rect 9690 -1442 10166 802
rect 12186 46 12392 1058
rect 12738 40 12944 1058
rect 13412 1054 13950 1058
rect 22971 1008 24060 1060
rect 14904 -1610 15172 796
rect 21882 -88 23078 -40
rect 21882 -216 21968 -88
rect 22960 -216 23078 -88
rect 21882 -248 23078 -216
rect 20054 -430 20494 -394
rect 20054 -506 20084 -430
rect 20462 -506 20494 -430
rect 20054 -510 20100 -506
rect 20446 -510 20494 -506
rect 20054 -540 20494 -510
rect 16228 -750 16616 -710
rect 16228 -1082 16268 -750
rect 16572 -1082 16616 -750
rect 16228 -1130 16616 -1082
rect 23638 -752 24060 1008
rect 23638 -1809 23696 -752
rect 944 -2052 1464 -1984
rect 20096 -1826 23696 -1809
rect 23998 -1826 24060 -752
rect 944 -2572 5348 -2052
rect 20096 -2231 24060 -1826
<< via3 >>
rect 3472 18152 7492 18612
rect 18164 18340 21510 18772
rect 11358 18188 11654 18322
rect 13410 18214 13932 18298
rect 2720 -238 3848 -90
rect 4368 -494 4880 -344
rect 8398 -1102 8632 -744
rect 21968 -216 22960 -88
rect 20084 -442 20462 -430
rect 20084 -504 20098 -442
rect 20098 -504 20442 -442
rect 20442 -504 20462 -442
rect 20084 -506 20462 -504
rect 20100 -510 20446 -506
rect 16268 -1082 16572 -750
<< metal4 >>
rect 13752 21330 24441 21898
rect 18057 18772 21688 18848
rect 3340 18612 7634 18650
rect 3340 18152 3472 18612
rect 7492 18152 7634 18612
rect 18057 18340 18164 18772
rect 21510 18340 21688 18772
rect 11282 18330 11684 18340
rect 10528 18322 11684 18330
rect 10528 18188 11358 18322
rect 11654 18188 11684 18322
rect 10528 18160 11684 18188
rect 13378 18298 14776 18314
rect 13378 18214 13410 18298
rect 13932 18214 14776 18298
rect 18057 18271 21688 18340
rect 13378 18182 14776 18214
rect 10528 18156 11604 18160
rect 3340 18086 7634 18152
rect 667 15985 1235 16520
rect 9294 16326 15970 16902
rect 23873 16320 24441 21330
rect 649 12201 1235 15985
rect 9306 14234 15754 14788
rect 667 -38 1235 12201
rect 9346 12142 15794 12696
rect 9274 10042 15722 10596
rect 9200 7982 16026 8526
rect 9170 5872 15996 6416
rect 11902 4332 15996 4346
rect 9170 3802 15996 4332
rect 9222 1670 16048 2214
rect 23771 -34 24339 2016
rect 667 -46 2952 -38
rect 22432 -40 24339 -34
rect 667 -90 3956 -46
rect 667 -238 2720 -90
rect 3848 -238 3956 -90
rect 667 -288 3956 -238
rect 21882 -88 24339 -40
rect 21882 -216 21968 -88
rect 22960 -216 24339 -88
rect 21882 -248 24339 -216
rect 22432 -260 24339 -248
rect 667 -302 2952 -288
rect 667 -2944 1235 -302
rect 4348 -344 4900 -326
rect 4348 -494 4368 -344
rect 4880 -410 4900 -344
rect 4880 -494 4904 -410
rect 4348 -512 4904 -494
rect 4366 -2044 4904 -512
rect 20054 -430 20494 -394
rect 20054 -506 20084 -430
rect 20462 -506 20494 -430
rect 20054 -510 20100 -506
rect 20446 -510 20494 -506
rect 20054 -540 20494 -510
rect 8366 -744 8664 -698
rect 8366 -1102 8398 -744
rect 8632 -1102 8664 -744
rect 8366 -1446 8664 -1102
rect 16224 -750 16610 -706
rect 16224 -1082 16268 -750
rect 16572 -1082 16610 -750
rect 16224 -1464 16610 -1082
rect 20062 -1924 20474 -540
rect 20630 -2014 20996 -2008
rect 23771 -2270 24339 -260
<< via4 >>
rect 3472 18152 7492 18612
rect 18164 18340 21510 18772
<< metal5 >>
rect 0 21211 11513 21801
rect 0 18625 590 21211
rect 18057 18772 25055 18861
rect 3340 18625 7634 18650
rect 0 18612 7634 18625
rect 0 18152 3472 18612
rect 7492 18152 7634 18612
rect 18057 18340 18164 18772
rect 21510 18340 25055 18772
rect 18057 18271 25055 18340
rect 0 18086 7634 18152
rect 0 18035 4377 18086
rect 0 14570 590 18035
rect 24465 16895 25055 18271
rect 9370 14854 16046 15430
rect 24465 14828 25083 16895
rect -8 14161 590 14570
rect -12 12853 590 14161
rect -12 12459 582 12853
rect 9294 12748 15742 13302
rect -12 11503 578 12459
rect -32 10235 578 11503
rect 9190 10658 15638 11212
rect -32 9379 558 10235
rect -32 798 572 9379
rect 9096 8568 15922 9112
rect 9054 6498 15880 7042
rect 9138 4408 15964 4952
rect 9138 2328 15964 2872
rect 24493 802 25083 14828
rect -32 194 2184 798
rect 22432 182 25083 802
rect 24493 -2270 25083 182
use capacitor_8  capacitor_8_0
timestamp 1698753667
transform 1 0 1274 0 1 182
box 0 -430 10546 2050
use capacitor_8  capacitor_8_1
timestamp 1698753667
transform -1 0 23730 0 1 194
box 0 -430 10546 2050
use capacitors_1  capacitors_1_0
timestamp 1698753667
transform 1 0 1295 0 1 14846
box -1291 -848 10655 2058
use capacitors_1  capacitors_1_1
timestamp 1698753667
transform -1 0 23807 0 1 14836
box -1291 -848 10655 2058
use capacitors_1  capacitors_1_2
timestamp 1698753667
transform 1 0 1265 0 1 12740
box -1291 -848 10655 2058
use capacitors_1  capacitors_1_3
timestamp 1698753667
transform 1 0 1269 0 1 10646
box -1291 -848 10655 2058
use capacitors_1  capacitors_1_4
timestamp 1698753667
transform -1 0 23799 0 1 12744
box -1291 -848 10655 2058
use capacitors_1  capacitors_1_5
timestamp 1698753667
transform -1 0 23775 0 1 10650
box -1291 -848 10655 2058
use capacitors_1  capacitors_1_6
timestamp 1698753667
transform 1 0 1261 0 1 8552
box -1291 -848 10655 2058
use capacitors_1  capacitors_1_7
timestamp 1698753667
transform 1 0 1251 0 1 6458
box -1291 -848 10655 2058
use capacitors_1  capacitors_1_8
timestamp 1698753667
transform 1 0 1251 0 1 4364
box -1291 -848 10655 2058
use capacitors_1  capacitors_1_9
timestamp 1698753667
transform 1 0 1263 0 1 2270
box -1291 -848 10655 2058
use capacitors_1  capacitors_1_10
timestamp 1698753667
transform -1 0 23705 0 1 2280
box -1291 -848 10655 2058
use capacitors_1  capacitors_1_11
timestamp 1698753667
transform -1 0 23727 0 1 4372
box -1291 -848 10655 2058
use capacitors_1  capacitors_1_12
timestamp 1698753667
transform -1 0 23791 0 1 6466
box -1291 -848 10655 2058
use capacitors_1  capacitors_1_13
timestamp 1698753667
transform -1 0 23831 0 1 8558
box -1291 -848 10655 2058
use clock  clock_1
timestamp 1698410772
transform 0 1 12960 -1 0 25486
box -410 -1832 6030 1274
use nmos_dnw3  nmos_dnw3_0
timestamp 1698467949
transform 1 0 12184 0 1 16340
box -424 892 1176 2258
use pmos_cp1  pmos_cp1_0
timestamp 1698464655
transform 1 0 12196 0 -1 182
box -14 -278 858 754
use sky130_fd_pr__cap_mim_m3_1_MH6KF8  sky130_fd_pr__cap_mim_m3_1_MH6KF8_0
timestamp 1698571947
transform -1 0 15980 0 1 -2156
box -1086 -940 1086 940
use sky130_fd_pr__cap_mim_m3_1_MH6KF8  sky130_fd_pr__cap_mim_m3_1_MH6KF8_1
timestamp 1698571947
transform 1 0 9038 0 1 -2176
box -1086 -940 1086 940
use sky130_fd_pr__cap_mim_m3_1_MH6KF8  sky130_fd_pr__cap_mim_m3_1_MH6KF8_2
timestamp 1698571947
transform 1 0 5164 0 1 -2412
box -1086 -940 1086 940
use sky130_fd_pr__cap_mim_m3_1_MH6KF8  sky130_fd_pr__cap_mim_m3_1_MH6KF8_3
timestamp 1698571947
transform -1 0 20174 0 1 -2456
box -1086 -940 1086 940
use sky130_fd_pr__cap_mim_m3_1_MH6KF8  sky130_fd_pr__cap_mim_m3_1_MH6KF8_4
timestamp 1698571947
transform -1 0 10140 0 1 18192
box -1086 -940 1086 940
use sky130_fd_pr__cap_mim_m3_1_MH6KF8  sky130_fd_pr__cap_mim_m3_1_MH6KF8_5
timestamp 1698571947
transform 1 0 15220 0 1 18184
box -1086 -940 1086 940
use sky130_fd_pr__nfet_01v8_NJGC8F  sky130_fd_pr__nfet_01v8_NJGC8F_0
timestamp 1698675553
transform 0 1 24518 -1 0 12713
box -3869 -130 3869 130
use sky130_fd_pr__nfet_01v8_NJGC8F  sky130_fd_pr__nfet_01v8_NJGC8F_1
timestamp 1698675553
transform 0 1 560 -1 0 4111
box -3869 -130 3869 130
use sky130_fd_pr__pfet_01v8_4RPJ49  sky130_fd_pr__pfet_01v8_4RPJ49_0
timestamp 1698675553
transform 0 1 24416 -1 0 4295
box -3905 -142 3905 142
use sky130_fd_pr__pfet_01v8_4RPJ49  sky130_fd_pr__pfet_01v8_4RPJ49_1
timestamp 1698675553
transform 0 1 670 -1 0 11955
box -3905 -142 3905 142
<< labels >>
rlabel metal3 12088 15446 12088 15446 1 input1
port 34 n
rlabel metal3 12964 15418 12964 15418 1 input2
port 35 n
rlabel metal4 964 12774 964 12774 1 vdd
port 1 n
rlabel metal5 24900 1146 24900 1146 1 gnd
port 64 n
rlabel metal2 12444 15904 12444 15904 1 in1
port 65 n
rlabel metal2 12576 11714 12576 11714 1 in3
port 66 n
rlabel metal2 12554 13796 12554 13796 1 in2
port 67 n
rlabel metal2 12598 9632 12598 9632 1 in4
port 68 n
rlabel metal2 12574 7544 12574 7544 1 in5
port 69 n
rlabel metal2 12526 5464 12526 5464 1 in6
port 70 n
rlabel metal2 12506 3382 12506 3382 1 in7
port 71 n
rlabel metal2 12554 1244 12554 1244 1 in8
port 73 n
<< end >>
