magic
tech sky130A
magscale 1 2
timestamp 1698771642
<< nmos >>
rect -927 -42 -897 42
rect -831 -42 -801 42
rect -735 -42 -705 42
rect -639 -42 -609 42
rect -543 -42 -513 42
rect -447 -42 -417 42
rect -351 -42 -321 42
rect -255 -42 -225 42
rect -159 -42 -129 42
rect -63 -42 -33 42
rect 33 -42 63 42
rect 129 -42 159 42
rect 225 -42 255 42
rect 321 -42 351 42
rect 417 -42 447 42
rect 513 -42 543 42
rect 609 -42 639 42
rect 705 -42 735 42
rect 801 -42 831 42
rect 897 -42 927 42
<< ndiff >>
rect -989 30 -927 42
rect -989 -30 -977 30
rect -943 -30 -927 30
rect -989 -42 -927 -30
rect -897 30 -831 42
rect -897 -30 -881 30
rect -847 -30 -831 30
rect -897 -42 -831 -30
rect -801 30 -735 42
rect -801 -30 -785 30
rect -751 -30 -735 30
rect -801 -42 -735 -30
rect -705 30 -639 42
rect -705 -30 -689 30
rect -655 -30 -639 30
rect -705 -42 -639 -30
rect -609 30 -543 42
rect -609 -30 -593 30
rect -559 -30 -543 30
rect -609 -42 -543 -30
rect -513 30 -447 42
rect -513 -30 -497 30
rect -463 -30 -447 30
rect -513 -42 -447 -30
rect -417 30 -351 42
rect -417 -30 -401 30
rect -367 -30 -351 30
rect -417 -42 -351 -30
rect -321 30 -255 42
rect -321 -30 -305 30
rect -271 -30 -255 30
rect -321 -42 -255 -30
rect -225 30 -159 42
rect -225 -30 -209 30
rect -175 -30 -159 30
rect -225 -42 -159 -30
rect -129 30 -63 42
rect -129 -30 -113 30
rect -79 -30 -63 30
rect -129 -42 -63 -30
rect -33 30 33 42
rect -33 -30 -17 30
rect 17 -30 33 30
rect -33 -42 33 -30
rect 63 30 129 42
rect 63 -30 79 30
rect 113 -30 129 30
rect 63 -42 129 -30
rect 159 30 225 42
rect 159 -30 175 30
rect 209 -30 225 30
rect 159 -42 225 -30
rect 255 30 321 42
rect 255 -30 271 30
rect 305 -30 321 30
rect 255 -42 321 -30
rect 351 30 417 42
rect 351 -30 367 30
rect 401 -30 417 30
rect 351 -42 417 -30
rect 447 30 513 42
rect 447 -30 463 30
rect 497 -30 513 30
rect 447 -42 513 -30
rect 543 30 609 42
rect 543 -30 559 30
rect 593 -30 609 30
rect 543 -42 609 -30
rect 639 30 705 42
rect 639 -30 655 30
rect 689 -30 705 30
rect 639 -42 705 -30
rect 735 30 801 42
rect 735 -30 751 30
rect 785 -30 801 30
rect 735 -42 801 -30
rect 831 30 897 42
rect 831 -30 847 30
rect 881 -30 897 30
rect 831 -42 897 -30
rect 927 30 989 42
rect 927 -30 943 30
rect 977 -30 989 30
rect 927 -42 989 -30
<< ndiffc >>
rect -977 -30 -943 30
rect -881 -30 -847 30
rect -785 -30 -751 30
rect -689 -30 -655 30
rect -593 -30 -559 30
rect -497 -30 -463 30
rect -401 -30 -367 30
rect -305 -30 -271 30
rect -209 -30 -175 30
rect -113 -30 -79 30
rect -17 -30 17 30
rect 79 -30 113 30
rect 175 -30 209 30
rect 271 -30 305 30
rect 367 -30 401 30
rect 463 -30 497 30
rect 559 -30 593 30
rect 655 -30 689 30
rect 751 -30 785 30
rect 847 -30 881 30
rect 943 -30 977 30
<< poly >>
rect -849 114 -783 130
rect -849 80 -833 114
rect -799 80 -783 114
rect -927 42 -897 68
rect -849 64 -783 80
rect -657 114 -591 130
rect -657 80 -641 114
rect -607 80 -591 114
rect -831 42 -801 64
rect -735 42 -705 68
rect -657 64 -591 80
rect -465 114 -399 130
rect -465 80 -449 114
rect -415 80 -399 114
rect -639 42 -609 64
rect -543 42 -513 68
rect -465 64 -399 80
rect -273 114 -207 130
rect -273 80 -257 114
rect -223 80 -207 114
rect -447 42 -417 64
rect -351 42 -321 68
rect -273 64 -207 80
rect -81 114 -15 130
rect -81 80 -65 114
rect -31 80 -15 114
rect -255 42 -225 64
rect -159 42 -129 68
rect -81 64 -15 80
rect 111 114 177 130
rect 111 80 127 114
rect 161 80 177 114
rect -63 42 -33 64
rect 33 42 63 68
rect 111 64 177 80
rect 303 114 369 130
rect 303 80 319 114
rect 353 80 369 114
rect 129 42 159 64
rect 225 42 255 68
rect 303 64 369 80
rect 495 114 561 130
rect 495 80 511 114
rect 545 80 561 114
rect 321 42 351 64
rect 417 42 447 68
rect 495 64 561 80
rect 687 114 753 130
rect 687 80 703 114
rect 737 80 753 114
rect 513 42 543 64
rect 609 42 639 68
rect 687 64 753 80
rect 879 114 945 130
rect 879 80 895 114
rect 929 80 945 114
rect 705 42 735 64
rect 801 42 831 68
rect 879 64 945 80
rect 897 42 927 64
rect -927 -64 -897 -42
rect -945 -80 -879 -64
rect -831 -68 -801 -42
rect -735 -64 -705 -42
rect -945 -114 -929 -80
rect -895 -114 -879 -80
rect -945 -130 -879 -114
rect -753 -80 -687 -64
rect -639 -68 -609 -42
rect -543 -64 -513 -42
rect -753 -114 -737 -80
rect -703 -114 -687 -80
rect -753 -130 -687 -114
rect -561 -80 -495 -64
rect -447 -68 -417 -42
rect -351 -64 -321 -42
rect -561 -114 -545 -80
rect -511 -114 -495 -80
rect -561 -130 -495 -114
rect -369 -80 -303 -64
rect -255 -68 -225 -42
rect -159 -64 -129 -42
rect -369 -114 -353 -80
rect -319 -114 -303 -80
rect -369 -130 -303 -114
rect -177 -80 -111 -64
rect -63 -68 -33 -42
rect 33 -64 63 -42
rect -177 -114 -161 -80
rect -127 -114 -111 -80
rect -177 -130 -111 -114
rect 15 -80 81 -64
rect 129 -68 159 -42
rect 225 -64 255 -42
rect 15 -114 31 -80
rect 65 -114 81 -80
rect 15 -130 81 -114
rect 207 -80 273 -64
rect 321 -68 351 -42
rect 417 -64 447 -42
rect 207 -114 223 -80
rect 257 -114 273 -80
rect 207 -130 273 -114
rect 399 -80 465 -64
rect 513 -68 543 -42
rect 609 -64 639 -42
rect 399 -114 415 -80
rect 449 -114 465 -80
rect 399 -130 465 -114
rect 591 -80 657 -64
rect 705 -68 735 -42
rect 801 -64 831 -42
rect 591 -114 607 -80
rect 641 -114 657 -80
rect 591 -130 657 -114
rect 783 -80 849 -64
rect 897 -68 927 -42
rect 783 -114 799 -80
rect 833 -114 849 -80
rect 783 -130 849 -114
<< polycont >>
rect -833 80 -799 114
rect -641 80 -607 114
rect -449 80 -415 114
rect -257 80 -223 114
rect -65 80 -31 114
rect 127 80 161 114
rect 319 80 353 114
rect 511 80 545 114
rect 703 80 737 114
rect 895 80 929 114
rect -929 -114 -895 -80
rect -737 -114 -703 -80
rect -545 -114 -511 -80
rect -353 -114 -319 -80
rect -161 -114 -127 -80
rect 31 -114 65 -80
rect 223 -114 257 -80
rect 415 -114 449 -80
rect 607 -114 641 -80
rect 799 -114 833 -80
<< locali >>
rect -849 80 -833 114
rect -799 80 -783 114
rect -657 80 -641 114
rect -607 80 -591 114
rect -465 80 -449 114
rect -415 80 -399 114
rect -273 80 -257 114
rect -223 80 -207 114
rect -81 80 -65 114
rect -31 80 -15 114
rect 111 80 127 114
rect 161 80 177 114
rect 303 80 319 114
rect 353 80 369 114
rect 495 80 511 114
rect 545 80 561 114
rect 687 80 703 114
rect 737 80 753 114
rect 879 80 895 114
rect 929 80 945 114
rect -977 30 -943 46
rect -977 -46 -943 -30
rect -881 30 -847 46
rect -881 -46 -847 -30
rect -785 30 -751 46
rect -785 -46 -751 -30
rect -689 30 -655 46
rect -689 -46 -655 -30
rect -593 30 -559 46
rect -593 -46 -559 -30
rect -497 30 -463 46
rect -497 -46 -463 -30
rect -401 30 -367 46
rect -401 -46 -367 -30
rect -305 30 -271 46
rect -305 -46 -271 -30
rect -209 30 -175 46
rect -209 -46 -175 -30
rect -113 30 -79 46
rect -113 -46 -79 -30
rect -17 30 17 46
rect -17 -46 17 -30
rect 79 30 113 46
rect 79 -46 113 -30
rect 175 30 209 46
rect 175 -46 209 -30
rect 271 30 305 46
rect 271 -46 305 -30
rect 367 30 401 46
rect 367 -46 401 -30
rect 463 30 497 46
rect 463 -46 497 -30
rect 559 30 593 46
rect 559 -46 593 -30
rect 655 30 689 46
rect 655 -46 689 -30
rect 751 30 785 46
rect 751 -46 785 -30
rect 847 30 881 46
rect 847 -46 881 -30
rect 943 30 977 46
rect 943 -46 977 -30
rect -945 -114 -929 -80
rect -895 -114 -879 -80
rect -753 -114 -737 -80
rect -703 -114 -687 -80
rect -561 -114 -545 -80
rect -511 -114 -495 -80
rect -369 -114 -353 -80
rect -319 -114 -303 -80
rect -177 -114 -161 -80
rect -127 -114 -111 -80
rect 15 -114 31 -80
rect 65 -114 81 -80
rect 207 -114 223 -80
rect 257 -114 273 -80
rect 399 -114 415 -80
rect 449 -114 465 -80
rect 591 -114 607 -80
rect 641 -114 657 -80
rect 783 -114 799 -80
rect 833 -114 849 -80
<< viali >>
rect -977 -30 -943 30
rect -881 -30 -847 30
rect -785 -30 -751 30
rect -689 -30 -655 30
rect -593 -30 -559 30
rect -497 -30 -463 30
rect -401 -30 -367 30
rect -305 -30 -271 30
rect -209 -30 -175 30
rect -113 -30 -79 30
rect -17 -30 17 30
rect 79 -30 113 30
rect 175 -30 209 30
rect 271 -30 305 30
rect 367 -30 401 30
rect 463 -30 497 30
rect 559 -30 593 30
rect 655 -30 689 30
rect 751 -30 785 30
rect 847 -30 881 30
rect 943 -30 977 30
<< metal1 >>
rect -983 30 -937 42
rect -983 -30 -977 30
rect -943 -30 -937 30
rect -983 -42 -937 -30
rect -887 30 -841 42
rect -887 -30 -881 30
rect -847 -30 -841 30
rect -887 -42 -841 -30
rect -791 30 -745 42
rect -791 -30 -785 30
rect -751 -30 -745 30
rect -791 -42 -745 -30
rect -695 30 -649 42
rect -695 -30 -689 30
rect -655 -30 -649 30
rect -695 -42 -649 -30
rect -599 30 -553 42
rect -599 -30 -593 30
rect -559 -30 -553 30
rect -599 -42 -553 -30
rect -503 30 -457 42
rect -503 -30 -497 30
rect -463 -30 -457 30
rect -503 -42 -457 -30
rect -407 30 -361 42
rect -407 -30 -401 30
rect -367 -30 -361 30
rect -407 -42 -361 -30
rect -311 30 -265 42
rect -311 -30 -305 30
rect -271 -30 -265 30
rect -311 -42 -265 -30
rect -215 30 -169 42
rect -215 -30 -209 30
rect -175 -30 -169 30
rect -215 -42 -169 -30
rect -119 30 -73 42
rect -119 -30 -113 30
rect -79 -30 -73 30
rect -119 -42 -73 -30
rect -23 30 23 42
rect -23 -30 -17 30
rect 17 -30 23 30
rect -23 -42 23 -30
rect 73 30 119 42
rect 73 -30 79 30
rect 113 -30 119 30
rect 73 -42 119 -30
rect 169 30 215 42
rect 169 -30 175 30
rect 209 -30 215 30
rect 169 -42 215 -30
rect 265 30 311 42
rect 265 -30 271 30
rect 305 -30 311 30
rect 265 -42 311 -30
rect 361 30 407 42
rect 361 -30 367 30
rect 401 -30 407 30
rect 361 -42 407 -30
rect 457 30 503 42
rect 457 -30 463 30
rect 497 -30 503 30
rect 457 -42 503 -30
rect 553 30 599 42
rect 553 -30 559 30
rect 593 -30 599 30
rect 553 -42 599 -30
rect 649 30 695 42
rect 649 -30 655 30
rect 689 -30 695 30
rect 649 -42 695 -30
rect 745 30 791 42
rect 745 -30 751 30
rect 785 -30 791 30
rect 745 -42 791 -30
rect 841 30 887 42
rect 841 -30 847 30
rect 881 -30 887 30
rect 841 -42 887 -30
rect 937 30 983 42
rect 937 -30 943 30
rect 977 -30 983 30
rect 937 -42 983 -30
<< properties >>
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 0.420 l 0.150 m 1 nf 20 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 0 botc 0 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 0 viasrc 100 viadrn 100 viagate 0 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
