magic
tech sky130A
magscale 1 2
timestamp 1698869963
<< metal2 >>
rect 22536 28901 23778 29141
rect 23538 28338 23778 28901
rect 69476 28867 70782 29107
rect 70542 28290 70782 28867
rect -1918 27158 1826 27230
rect 21640 27154 25190 27212
rect 45120 27134 48796 27218
rect 68590 27124 72170 27192
rect -1912 25076 1832 25148
rect 21632 25068 25182 25126
rect 45104 25044 48780 25128
rect 68580 25032 72160 25100
rect -1926 22992 1818 23064
rect 21592 22974 25244 23036
rect 45112 22946 48788 23030
rect 68584 22934 72164 23002
rect -1984 20896 1760 20968
rect 21614 20884 25266 20946
rect 45044 20862 48720 20946
rect 68570 20850 72150 20918
rect -2006 18798 1738 18870
rect 21626 18784 25278 18846
rect 45030 18772 48706 18856
rect 68590 18756 72170 18824
rect -2006 16716 1738 16788
rect 21692 16690 25268 16760
rect 45022 16674 48698 16758
rect 68670 16674 72250 16742
rect -1992 14626 1752 14698
rect 21710 14600 25286 14670
rect 45000 14568 48676 14652
rect 68656 14566 72236 14634
rect -1998 12514 1746 12586
rect 21710 12518 25286 12588
rect 45030 12484 48706 12568
rect 68676 12434 72226 12554
rect -130 10857 110 11462
rect -982 10617 110 10857
rect 46894 10831 47134 11394
rect 46178 10591 47134 10831
<< metal3 >>
rect -1234 975 390 1367
rect 21128 987 25434 1379
rect 43352 941 48538 1333
rect 68120 963 72286 1355
<< metal4 >>
rect -24265 28249 -23567 28279
rect -24265 27695 -12961 28249
rect -24265 26161 -23567 27695
rect 83365 27651 94515 28205
rect -24265 25607 -12413 26161
rect 93961 26117 94515 27651
rect -24265 24093 -23567 25607
rect 82883 25563 94515 26117
rect -24265 23539 -12515 24093
rect 93961 24049 94515 25563
rect -24265 21999 -23567 23539
rect 83095 23495 94515 24049
rect -24265 21445 -12433 21999
rect 93961 21955 94515 23495
rect -24265 19883 -23567 21445
rect 83265 21401 94515 21955
rect -24265 19329 -12403 19883
rect 93961 19839 94515 21401
rect -24265 17829 -23567 19329
rect 83115 19285 94515 19839
rect -24265 17275 -12341 17829
rect 93961 17785 94515 19285
rect -24265 15761 -23567 17275
rect 82933 17231 94515 17785
rect -24265 15724 -21280 15761
rect -13716 15738 -12707 15761
rect -15656 15724 -12707 15738
rect -24265 15207 -12707 15724
rect 93961 15717 94515 17231
rect 85904 15694 85906 15698
rect 82903 15662 85906 15694
rect 91566 15662 94515 15717
rect -24265 13659 -23567 15207
rect 82903 15163 94515 15662
rect -24265 13105 -12595 13659
rect 93961 13615 94515 15163
rect -24265 6682 -23567 13105
rect 83145 13061 94515 13615
rect -24284 6031 -15911 6682
rect -24265 2170 -23567 6031
rect -24265 1472 -13560 2170
rect -1397 1450 696 2148
rect 20917 1444 25977 2142
rect 93961 2120 94515 13061
rect 43493 1416 49395 2114
rect 67341 1420 73163 2118
rect 82277 1422 94539 2120
<< metal5 >>
rect -25261 26777 -24543 26811
rect -25261 26223 -12759 26777
rect -25261 24681 -24543 26223
rect 92084 26189 95040 26761
rect -25261 24127 -12909 24681
rect 94468 24637 95040 26189
rect -25261 22607 -24543 24127
rect 83297 24083 95040 24637
rect -25261 22053 -12257 22607
rect 94468 22563 95040 24083
rect -25261 20527 -24543 22053
rect 83105 22009 95040 22563
rect -25261 19973 -12289 20527
rect 94468 20483 95040 22009
rect -25261 18445 -24543 19973
rect 82945 19929 95040 20483
rect -25261 17891 -12257 18445
rect 94468 18401 95040 19929
rect -25261 16371 -24543 17891
rect 83025 17847 95113 18401
rect -25261 15817 -12385 16371
rect 94468 16327 95040 17847
rect -25261 14255 -24543 15817
rect 83125 15773 95040 16327
rect -25261 13701 -12343 14255
rect 94468 14211 95040 15773
rect -25261 12201 -24543 13701
rect 82743 13657 95040 14211
rect -25261 11647 -12835 12201
rect 94468 12157 95040 13657
rect -25261 894 -24543 11647
rect 83105 11603 95081 12157
rect -25261 176 -19513 894
rect -889 156 1175 835
rect 21709 150 26985 868
rect 44363 122 48034 801
rect 68133 126 73193 844
rect 94468 805 95040 11603
rect 91983 126 95043 805
use cp2_buffer1  cp2_buffer1_0
timestamp 1698849032
transform 1 0 -27092 0 1 1943
box 3710 -1785 26750 28454
use cp2_buffer1  cp2_buffer1_1
timestamp 1698849032
transform 1 0 19930 0 1 1917
box 3710 -1785 26750 28454
use cp2_buffer1  cp2_buffer1_2
timestamp 1698849032
transform 1 0 66898 0 1 1893
box 3710 -1785 26750 28454
use cp2_buffer2  cp2_buffer2_0
timestamp 1698869963
transform 1 0 -28016 0 1 1923
box 28006 -1775 51269 29658
use cp2_buffer2  cp2_buffer2_1
timestamp 1698869963
transform 1 0 18930 0 1 1889
box 28006 -1775 51269 29658
<< end >>
