magic
tech sky130A
magscale 1 2
timestamp 1699075837
<< nwell >>
rect -114 1010 368 1466
rect -114 994 238 1010
rect -114 990 -80 994
<< psubdiff >>
rect 34 744 148 766
rect 34 646 64 744
rect 122 646 148 744
rect 34 616 148 646
<< nsubdiff >>
rect -28 1376 68 1418
rect -28 1204 -6 1376
rect 48 1204 68 1376
rect -28 1164 68 1204
<< psubdiffcont >>
rect 64 646 122 744
<< nsubdiffcont >>
rect -6 1204 48 1376
<< poly >>
rect 744 114 2590 156
rect 740 90 2590 114
rect 740 20 2598 90
rect 6494 68 7422 112
rect 740 -8 770 20
rect 932 -12 962 20
rect 1124 -6 1154 20
rect 1316 -8 1346 20
rect 1508 -12 1538 20
rect 1700 -18 1730 20
rect 1892 -8 1922 20
rect 1892 -16 1922 -10
rect 2084 -16 2114 20
rect 2276 -20 2306 20
rect 2468 -10 2498 20
rect 3022 -34 3052 -10
rect 3214 -34 3244 -10
rect 3406 -34 3436 12
rect 3598 -34 3628 8
rect 3790 -34 3820 4
rect 3982 -34 4012 0
rect 4174 -34 4204 10
rect 4366 -34 4396 4
rect 4558 -34 4588 14
rect 4750 -34 4780 2
rect 2858 -174 4840 -34
rect 5452 -56 5482 20
rect 5644 -56 5674 16
rect 5836 -56 5866 20
rect 6028 -56 6058 16
rect 6220 -56 6250 16
rect 6480 4 7422 68
rect 6480 -30 6510 4
rect 6672 -32 6702 4
rect 6864 -34 6894 4
rect 7056 -34 7086 4
rect 7248 -38 7278 4
rect 5270 -86 6302 -56
rect 5270 -124 6278 -86
<< locali >>
rect -28 1376 68 1418
rect -28 1204 -6 1376
rect 48 1204 68 1376
rect -28 1164 68 1204
rect 34 744 148 766
rect 34 646 64 744
rect 122 646 148 744
rect 34 616 148 646
rect 744 486 2702 522
rect 744 364 2590 486
rect 744 246 896 364
rect 742 184 896 246
rect 2462 184 2590 364
rect 742 90 2590 184
rect 6492 442 7386 524
rect 6492 148 6554 442
rect 7308 148 7386 442
rect 6492 112 7386 148
rect 742 88 2598 90
rect 792 20 2598 88
rect 6492 52 7422 112
rect 6494 4 7422 52
rect 2858 -134 4840 -42
rect 2858 -182 2922 -134
rect 2872 -384 2922 -182
rect 4672 -182 4840 -134
rect 5270 -140 6302 -56
rect 4672 -384 4832 -182
rect 2872 -416 4832 -384
rect 5270 -382 5304 -140
rect 6250 -382 6302 -140
rect 5270 -402 6302 -382
<< viali >>
rect -6 1204 48 1376
rect 64 646 122 744
rect 896 184 2462 364
rect 6554 148 7308 442
rect 2922 -384 4672 -134
rect 5304 -382 6250 -140
<< metal1 >>
rect -338 2046 362 2047
rect -534 1944 362 2046
rect -534 1820 536 1944
rect -534 1584 496 1820
rect -534 1472 268 1584
rect -534 1470 -102 1472
rect -466 1319 -432 1470
rect -248 1315 -214 1470
rect -28 1376 66 1472
rect -28 1204 -6 1376
rect 48 1204 66 1376
rect -28 1164 66 1204
rect -94 1000 240 1006
rect -94 990 -68 1000
rect -96 948 -68 990
rect -94 940 -68 948
rect 192 940 240 1000
rect -94 932 240 940
rect 7200 930 7656 948
rect 7200 870 7216 930
rect 7108 850 7216 870
rect 7608 850 7656 930
rect 7108 838 7656 850
rect -466 796 -432 834
rect -248 796 -214 834
rect -530 548 -58 796
rect 34 766 146 768
rect 34 744 148 766
rect 34 646 64 744
rect 122 646 148 744
rect 34 616 148 646
rect 34 548 146 616
rect -530 522 438 548
rect 6338 534 7541 568
rect 5290 530 7541 534
rect -531 488 2702 522
rect 2824 506 4846 514
rect 2824 488 4880 506
rect -531 474 1168 488
rect 2588 474 2598 484
rect -531 364 2598 474
rect -531 184 896 364
rect 2462 184 2598 364
rect -531 88 2598 184
rect 2836 140 4880 488
rect 782 86 2598 88
rect 2834 80 4880 140
rect 3274 -2 4880 80
rect 5282 442 7541 530
rect 5282 148 6554 442
rect 7308 148 7541 442
rect 5282 3 7541 148
rect 3274 -4 3362 -2
rect 5282 -8 6338 3
rect 602 -334 2650 -60
rect 2810 -134 4832 -68
rect 2810 -384 2922 -134
rect 4672 -384 4832 -134
rect 2810 -430 4832 -384
rect 5270 -140 6302 -56
rect 5270 -382 5304 -140
rect 6250 -382 6302 -140
rect 6370 -278 7460 -54
rect 5270 -402 6302 -382
<< via1 >>
rect -68 940 192 1000
rect 7216 850 7608 930
<< metal2 >>
rect 340 1084 536 1086
rect 164 1082 536 1084
rect -739 1036 9792 1082
rect -738 930 -694 1036
rect 7406 1030 9792 1036
rect -94 1000 240 1006
rect -94 990 -68 1000
rect -96 948 -68 990
rect -94 940 -68 948
rect 192 940 240 1000
rect -94 932 240 940
rect 7200 930 7634 948
rect 7200 850 7216 930
rect 7608 850 7634 930
rect 7200 838 7634 850
<< via2 >>
rect 7216 850 7608 930
<< metal3 >>
rect 7758 966 9428 1828
rect 7200 930 7634 948
rect 7200 850 7216 930
rect 7608 850 7634 930
rect 7200 838 7634 850
rect 7758 720 9807 966
rect 7758 166 9428 720
<< via3 >>
rect 7216 850 7608 930
<< mimcap >>
rect 7800 932 9394 1798
rect 7800 839 7999 932
rect 7800 762 7838 839
rect 8118 762 9394 932
rect 7800 200 9394 762
<< mimcapcontact >>
rect 7999 839 8118 932
rect 7838 762 8118 839
<< metal4 >>
rect 7999 953 8144 954
rect 7758 950 8144 953
rect 7200 932 8144 950
rect 7200 930 7999 932
rect 7200 850 7216 930
rect 7608 850 7999 930
rect 7200 839 7999 850
rect 7200 838 7838 839
rect 7758 762 7838 838
rect 8118 762 8144 932
rect 7758 726 8144 762
use buffer_and_gate  buffer_and_gate_0
timestamp 1698998396
transform 1 0 84 0 1 30
box -116 -30 7470 2020
use buffer_digital  buffer_digital_0
timestamp 1699074083
transform 1 0 -464 0 1 800
box -274 -74 412 576
use sky130_fd_pr__nfet_01v8_9LGCGE  sky130_fd_pr__nfet_01v8_9LGCGE_0
timestamp 1699075837
transform 1 0 3853 0 1 38
box -989 -130 989 130
use sky130_fd_pr__nfet_01v8_NJGC45  sky130_fd_pr__nfet_01v8_NJGC45_0
timestamp 1698837560
transform 1 0 5803 0 1 26
box -509 -130 509 130
use sky130_fd_pr__pfet_01v8_4ZKXAA  sky130_fd_pr__pfet_01v8_4ZKXAA_0
timestamp 1698837886
transform 1 0 6927 0 1 -88
box -545 -142 545 142
use sky130_fd_pr__pfet_01v8_49FP49  sky130_fd_pr__pfet_01v8_49FP49_0
timestamp 1698771642
transform 1 0 1667 0 1 -70
box -1025 -142 1025 142
<< end >>
