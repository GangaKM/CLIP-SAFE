magic
tech sky130A
magscale 1 2
timestamp 1698756166
<< nwell >>
rect 23810 -2372 24396 -1994
rect 29962 -2380 30562 -1916
rect 47806 -2372 48466 -1994
rect 54248 -2382 54840 -2002
rect 73810 -2472 74456 -2096
rect 80100 -2106 80768 -2100
rect 80100 -2482 80834 -2106
rect 99805 -2272 100560 -1895
rect 106201 -2282 106834 -1902
<< nmos >>
rect 47904 -2524 47934 -2440
rect 48122 -2524 48152 -2440
rect 54492 -2534 54522 -2450
rect 54710 -2534 54740 -2450
rect 99904 -2424 99934 -2340
rect 100122 -2424 100152 -2340
rect 106492 -2434 106522 -2350
rect 106710 -2434 106740 -2350
rect 73904 -2624 73934 -2540
rect 74122 -2624 74152 -2540
rect 80492 -2634 80522 -2550
rect 80710 -2634 80740 -2550
<< pmos >>
rect 47904 -2310 47934 -2058
rect 48122 -2310 48152 -2058
rect 54492 -2320 54522 -2068
rect 54710 -2320 54740 -2068
rect 73904 -2410 73934 -2158
rect 74122 -2410 74152 -2158
rect 80492 -2420 80522 -2168
rect 80710 -2420 80740 -2168
rect 99904 -2210 99934 -1958
rect 100122 -2210 100152 -1958
rect 106492 -2220 106522 -1968
rect 106710 -2220 106740 -1968
<< ndiff >>
rect 47846 -2452 47904 -2440
rect 47846 -2512 47858 -2452
rect 47892 -2512 47904 -2452
rect 47846 -2524 47904 -2512
rect 47934 -2452 47992 -2440
rect 47934 -2512 47946 -2452
rect 47980 -2512 47992 -2452
rect 47934 -2524 47992 -2512
rect 48064 -2452 48122 -2440
rect 48064 -2512 48076 -2452
rect 48110 -2512 48122 -2452
rect 48064 -2524 48122 -2512
rect 48152 -2452 48210 -2440
rect 48152 -2512 48164 -2452
rect 48198 -2512 48210 -2452
rect 48152 -2524 48210 -2512
rect 54434 -2462 54492 -2450
rect 54434 -2522 54446 -2462
rect 54480 -2522 54492 -2462
rect 54434 -2534 54492 -2522
rect 54522 -2462 54580 -2450
rect 54522 -2522 54534 -2462
rect 54568 -2522 54580 -2462
rect 54522 -2534 54580 -2522
rect 54652 -2462 54710 -2450
rect 54652 -2522 54664 -2462
rect 54698 -2522 54710 -2462
rect 54652 -2534 54710 -2522
rect 54740 -2462 54798 -2450
rect 54740 -2522 54752 -2462
rect 54786 -2522 54798 -2462
rect 99846 -2352 99904 -2340
rect 99846 -2412 99858 -2352
rect 99892 -2412 99904 -2352
rect 54740 -2534 54798 -2522
rect 99846 -2424 99904 -2412
rect 99934 -2352 99992 -2340
rect 99934 -2412 99946 -2352
rect 99980 -2412 99992 -2352
rect 99934 -2424 99992 -2412
rect 100064 -2352 100122 -2340
rect 100064 -2412 100076 -2352
rect 100110 -2412 100122 -2352
rect 100064 -2424 100122 -2412
rect 100152 -2352 100210 -2340
rect 100152 -2412 100164 -2352
rect 100198 -2412 100210 -2352
rect 100152 -2424 100210 -2412
rect 106434 -2362 106492 -2350
rect 106434 -2422 106446 -2362
rect 106480 -2422 106492 -2362
rect 106434 -2434 106492 -2422
rect 106522 -2362 106580 -2350
rect 106522 -2422 106534 -2362
rect 106568 -2422 106580 -2362
rect 106522 -2434 106580 -2422
rect 106652 -2362 106710 -2350
rect 106652 -2422 106664 -2362
rect 106698 -2422 106710 -2362
rect 106652 -2434 106710 -2422
rect 106740 -2362 106798 -2350
rect 106740 -2422 106752 -2362
rect 106786 -2422 106798 -2362
rect 106740 -2434 106798 -2422
rect 73846 -2552 73904 -2540
rect 73846 -2612 73858 -2552
rect 73892 -2612 73904 -2552
rect 73846 -2624 73904 -2612
rect 73934 -2552 73992 -2540
rect 73934 -2612 73946 -2552
rect 73980 -2612 73992 -2552
rect 73934 -2624 73992 -2612
rect 74064 -2552 74122 -2540
rect 74064 -2612 74076 -2552
rect 74110 -2612 74122 -2552
rect 74064 -2624 74122 -2612
rect 74152 -2552 74210 -2540
rect 74152 -2612 74164 -2552
rect 74198 -2612 74210 -2552
rect 74152 -2624 74210 -2612
rect 80434 -2562 80492 -2550
rect 80434 -2622 80446 -2562
rect 80480 -2622 80492 -2562
rect 80434 -2634 80492 -2622
rect 80522 -2562 80580 -2550
rect 80522 -2622 80534 -2562
rect 80568 -2622 80580 -2562
rect 80522 -2634 80580 -2622
rect 80652 -2562 80710 -2550
rect 80652 -2622 80664 -2562
rect 80698 -2622 80710 -2562
rect 80652 -2634 80710 -2622
rect 80740 -2562 80798 -2550
rect 80740 -2622 80752 -2562
rect 80786 -2622 80798 -2562
rect 80740 -2634 80798 -2622
<< pdiff >>
rect 99846 -1970 99904 -1958
rect 47846 -2070 47904 -2058
rect 47846 -2298 47858 -2070
rect 47892 -2298 47904 -2070
rect 47846 -2310 47904 -2298
rect 47934 -2070 47992 -2058
rect 47934 -2298 47946 -2070
rect 47980 -2298 47992 -2070
rect 47934 -2310 47992 -2298
rect 48064 -2070 48122 -2058
rect 48064 -2298 48076 -2070
rect 48110 -2298 48122 -2070
rect 48064 -2310 48122 -2298
rect 48152 -2070 48210 -2058
rect 48152 -2298 48164 -2070
rect 48198 -2298 48210 -2070
rect 54434 -2080 54492 -2068
rect 48152 -2310 48210 -2298
rect 54434 -2308 54446 -2080
rect 54480 -2308 54492 -2080
rect 54434 -2320 54492 -2308
rect 54522 -2080 54580 -2068
rect 54522 -2308 54534 -2080
rect 54568 -2308 54580 -2080
rect 54522 -2320 54580 -2308
rect 54652 -2080 54710 -2068
rect 54652 -2308 54664 -2080
rect 54698 -2308 54710 -2080
rect 54652 -2320 54710 -2308
rect 54740 -2080 54798 -2068
rect 54740 -2308 54752 -2080
rect 54786 -2308 54798 -2080
rect 54740 -2320 54798 -2308
rect 73846 -2170 73904 -2158
rect 73846 -2398 73858 -2170
rect 73892 -2398 73904 -2170
rect 73846 -2410 73904 -2398
rect 73934 -2170 73992 -2158
rect 73934 -2398 73946 -2170
rect 73980 -2398 73992 -2170
rect 73934 -2410 73992 -2398
rect 74064 -2170 74122 -2158
rect 74064 -2398 74076 -2170
rect 74110 -2398 74122 -2170
rect 74064 -2410 74122 -2398
rect 74152 -2170 74210 -2158
rect 74152 -2398 74164 -2170
rect 74198 -2398 74210 -2170
rect 80434 -2180 80492 -2168
rect 74152 -2410 74210 -2398
rect 80434 -2408 80446 -2180
rect 80480 -2408 80492 -2180
rect 80434 -2420 80492 -2408
rect 80522 -2180 80580 -2168
rect 80522 -2408 80534 -2180
rect 80568 -2408 80580 -2180
rect 80522 -2420 80580 -2408
rect 80652 -2180 80710 -2168
rect 80652 -2408 80664 -2180
rect 80698 -2408 80710 -2180
rect 80652 -2420 80710 -2408
rect 80740 -2180 80798 -2168
rect 80740 -2408 80752 -2180
rect 80786 -2408 80798 -2180
rect 99846 -2198 99858 -1970
rect 99892 -2198 99904 -1970
rect 99846 -2210 99904 -2198
rect 99934 -1970 99992 -1958
rect 99934 -2198 99946 -1970
rect 99980 -2198 99992 -1970
rect 99934 -2210 99992 -2198
rect 100064 -1970 100122 -1958
rect 100064 -2198 100076 -1970
rect 100110 -2198 100122 -1970
rect 100064 -2210 100122 -2198
rect 100152 -1970 100210 -1958
rect 100152 -2198 100164 -1970
rect 100198 -2198 100210 -1970
rect 106434 -1980 106492 -1968
rect 100152 -2210 100210 -2198
rect 106434 -2208 106446 -1980
rect 106480 -2208 106492 -1980
rect 106434 -2220 106492 -2208
rect 106522 -1980 106580 -1968
rect 106522 -2208 106534 -1980
rect 106568 -2208 106580 -1980
rect 106522 -2220 106580 -2208
rect 106652 -1980 106710 -1968
rect 106652 -2208 106664 -1980
rect 106698 -2208 106710 -1980
rect 106652 -2220 106710 -2208
rect 106740 -1980 106798 -1968
rect 106740 -2208 106752 -1980
rect 106786 -2208 106798 -1980
rect 106740 -2220 106798 -2208
rect 80740 -2420 80798 -2408
<< ndiffc >>
rect 47858 -2512 47892 -2452
rect 47946 -2512 47980 -2452
rect 48076 -2512 48110 -2452
rect 48164 -2512 48198 -2452
rect 54446 -2522 54480 -2462
rect 54534 -2522 54568 -2462
rect 54664 -2522 54698 -2462
rect 54752 -2522 54786 -2462
rect 99858 -2412 99892 -2352
rect 99946 -2412 99980 -2352
rect 100076 -2412 100110 -2352
rect 100164 -2412 100198 -2352
rect 106446 -2422 106480 -2362
rect 106534 -2422 106568 -2362
rect 106664 -2422 106698 -2362
rect 106752 -2422 106786 -2362
rect 73858 -2612 73892 -2552
rect 73946 -2612 73980 -2552
rect 74076 -2612 74110 -2552
rect 74164 -2612 74198 -2552
rect 80446 -2622 80480 -2562
rect 80534 -2622 80568 -2562
rect 80664 -2622 80698 -2562
rect 80752 -2622 80786 -2562
<< pdiffc >>
rect 47858 -2298 47892 -2070
rect 47946 -2298 47980 -2070
rect 48076 -2298 48110 -2070
rect 48164 -2298 48198 -2070
rect 54446 -2308 54480 -2080
rect 54534 -2308 54568 -2080
rect 54664 -2308 54698 -2080
rect 54752 -2308 54786 -2080
rect 73858 -2398 73892 -2170
rect 73946 -2398 73980 -2170
rect 74076 -2398 74110 -2170
rect 74164 -2398 74198 -2170
rect 80446 -2408 80480 -2180
rect 80534 -2408 80568 -2180
rect 80664 -2408 80698 -2180
rect 80752 -2408 80786 -2180
rect 99858 -2198 99892 -1970
rect 99946 -2198 99980 -1970
rect 100076 -2198 100110 -1970
rect 100164 -2198 100198 -1970
rect 106446 -2208 106480 -1980
rect 106534 -2208 106568 -1980
rect 106664 -2208 106698 -1980
rect 106752 -2208 106786 -1980
<< nsubdiff >>
rect 29998 -2156 30090 -2126
rect 24264 -2182 24350 -2158
rect 24264 -2216 24288 -2182
rect 24324 -2216 24350 -2182
rect 29998 -2192 30024 -2156
rect 30062 -2192 30090 -2156
rect 29998 -2216 30090 -2192
rect 24264 -2244 24350 -2216
rect 48292 -2164 48394 -2130
rect 48292 -2200 48320 -2164
rect 48362 -2200 48394 -2164
rect 48292 -2226 48394 -2200
rect 54286 -2184 54358 -2158
rect 54286 -2218 54304 -2184
rect 54340 -2218 54358 -2184
rect 54286 -2246 54358 -2218
rect 74292 -2278 74374 -2236
rect 74292 -2318 74312 -2278
rect 74350 -2318 74374 -2278
rect 74292 -2344 74374 -2318
rect 80179 -2277 80303 -2242
rect 80179 -2337 80211 -2277
rect 80267 -2337 80303 -2277
rect 80179 -2371 80303 -2337
rect 100342 -2070 100457 -2036
rect 100342 -2122 100370 -2070
rect 100424 -2122 100457 -2070
rect 100342 -2152 100457 -2122
rect 106247 -2097 106346 -2065
rect 106247 -2139 106271 -2097
rect 106313 -2139 106346 -2097
rect 106247 -2161 106346 -2139
<< nsubdiffcont >>
rect 24288 -2216 24324 -2182
rect 30024 -2192 30062 -2156
rect 48320 -2200 48362 -2164
rect 54304 -2218 54340 -2184
rect 74312 -2318 74350 -2278
rect 80211 -2337 80267 -2277
rect 100370 -2122 100424 -2070
rect 106271 -2139 106313 -2097
<< poly >>
rect 99904 -1958 99934 -1932
rect 100122 -1958 100152 -1932
rect 47904 -2058 47934 -2032
rect 48122 -2058 48152 -2032
rect 47258 -2158 47674 -2116
rect 47258 -2618 47332 -2158
rect 47596 -2368 47674 -2158
rect 54492 -2068 54522 -2042
rect 54710 -2068 54740 -2042
rect 47904 -2368 47934 -2310
rect 48122 -2348 48152 -2310
rect 73904 -2158 73934 -2132
rect 74122 -2158 74152 -2132
rect 47596 -2400 47934 -2368
rect 47596 -2618 47674 -2400
rect 47904 -2440 47934 -2400
rect 47976 -2358 48152 -2348
rect 47976 -2394 48000 -2358
rect 48102 -2394 48152 -2358
rect 47976 -2404 48152 -2394
rect 48122 -2440 48152 -2404
rect 54174 -2376 54406 -2360
rect 54174 -2416 54192 -2376
rect 54386 -2378 54406 -2376
rect 54492 -2378 54522 -2320
rect 54710 -2358 54740 -2320
rect 54386 -2410 54522 -2378
rect 54386 -2416 54406 -2410
rect 54174 -2432 54406 -2416
rect 54492 -2450 54522 -2410
rect 54564 -2368 54740 -2358
rect 54564 -2404 54588 -2368
rect 54690 -2404 54740 -2368
rect 54564 -2414 54740 -2404
rect 80492 -2168 80522 -2142
rect 80710 -2168 80740 -2142
rect 54710 -2450 54740 -2414
rect 47904 -2550 47934 -2524
rect 48122 -2550 48152 -2524
rect 73586 -2466 73818 -2450
rect 73586 -2506 73604 -2466
rect 73798 -2468 73818 -2466
rect 73904 -2468 73934 -2410
rect 74122 -2448 74152 -2410
rect 106492 -1968 106522 -1942
rect 106710 -1968 106740 -1942
rect 99586 -2266 99818 -2250
rect 99586 -2306 99604 -2266
rect 99798 -2268 99818 -2266
rect 99904 -2268 99934 -2210
rect 100122 -2248 100152 -2210
rect 99798 -2300 99934 -2268
rect 99798 -2306 99818 -2300
rect 99586 -2322 99818 -2306
rect 99904 -2340 99934 -2300
rect 99976 -2258 100152 -2248
rect 99976 -2294 100000 -2258
rect 100102 -2294 100152 -2258
rect 99976 -2304 100152 -2294
rect 100122 -2340 100152 -2304
rect 106174 -2276 106406 -2260
rect 106174 -2316 106192 -2276
rect 106386 -2278 106406 -2276
rect 106492 -2278 106522 -2220
rect 106710 -2258 106740 -2220
rect 106386 -2310 106522 -2278
rect 106386 -2316 106406 -2310
rect 106174 -2332 106406 -2316
rect 73798 -2500 73934 -2468
rect 73798 -2506 73818 -2500
rect 73586 -2522 73818 -2506
rect 54492 -2560 54522 -2534
rect 54710 -2560 54740 -2534
rect 73904 -2540 73934 -2500
rect 73976 -2458 74152 -2448
rect 73976 -2494 74000 -2458
rect 74102 -2494 74152 -2458
rect 73976 -2504 74152 -2494
rect 74122 -2540 74152 -2504
rect 80174 -2476 80406 -2460
rect 80174 -2516 80192 -2476
rect 80386 -2478 80406 -2476
rect 80492 -2478 80522 -2420
rect 80710 -2458 80740 -2420
rect 106492 -2350 106522 -2310
rect 106564 -2268 106740 -2258
rect 106564 -2304 106588 -2268
rect 106690 -2304 106740 -2268
rect 106564 -2314 106740 -2304
rect 106710 -2350 106740 -2314
rect 99904 -2450 99934 -2424
rect 100122 -2450 100152 -2424
rect 80386 -2510 80522 -2478
rect 80386 -2516 80406 -2510
rect 80174 -2532 80406 -2516
rect 47258 -2656 47674 -2618
rect 80492 -2550 80522 -2510
rect 80564 -2468 80740 -2458
rect 106492 -2460 106522 -2434
rect 106710 -2460 106740 -2434
rect 80564 -2504 80588 -2468
rect 80690 -2504 80740 -2468
rect 80564 -2514 80740 -2504
rect 80710 -2550 80740 -2514
rect 73904 -2650 73934 -2624
rect 74122 -2650 74152 -2624
rect 80492 -2660 80522 -2634
rect 80710 -2660 80740 -2634
<< polycont >>
rect 47332 -2618 47596 -2158
rect 48000 -2394 48102 -2358
rect 54192 -2416 54386 -2376
rect 54588 -2404 54690 -2368
rect 73604 -2506 73798 -2466
rect 99604 -2306 99798 -2266
rect 100000 -2294 100102 -2258
rect 106192 -2316 106386 -2276
rect 74000 -2494 74102 -2458
rect 80192 -2516 80386 -2476
rect 106588 -2304 106690 -2268
rect 80588 -2504 80690 -2468
<< locali >>
rect 99858 -1970 99892 -1954
rect 47858 -2070 47892 -2054
rect 29998 -2156 30090 -2126
rect 24264 -2182 24350 -2158
rect 24264 -2216 24288 -2182
rect 24324 -2216 24350 -2182
rect 29998 -2192 30024 -2156
rect 30062 -2192 30090 -2156
rect 29998 -2216 30090 -2192
rect 47258 -2158 47674 -2116
rect 24264 -2244 24350 -2216
rect 47258 -2618 47332 -2158
rect 47596 -2618 47674 -2158
rect 47858 -2314 47892 -2298
rect 47946 -2070 47980 -2054
rect 47946 -2314 47980 -2298
rect 48076 -2070 48110 -2054
rect 48076 -2314 48110 -2298
rect 48164 -2070 48198 -2054
rect 54446 -2080 54480 -2064
rect 48292 -2164 48394 -2130
rect 48292 -2200 48320 -2164
rect 48362 -2200 48394 -2164
rect 48292 -2226 48394 -2200
rect 54286 -2184 54358 -2158
rect 54286 -2218 54304 -2184
rect 54340 -2218 54358 -2184
rect 54286 -2246 54358 -2218
rect 48164 -2314 48198 -2298
rect 54446 -2324 54480 -2308
rect 54534 -2080 54568 -2064
rect 54534 -2324 54568 -2308
rect 54664 -2080 54698 -2064
rect 54664 -2324 54698 -2308
rect 54752 -2080 54786 -2064
rect 54752 -2324 54786 -2308
rect 73858 -2170 73892 -2154
rect 47976 -2358 48134 -2348
rect 47976 -2394 48000 -2358
rect 48102 -2394 48134 -2358
rect 47976 -2402 48134 -2394
rect 54174 -2376 54406 -2360
rect 54174 -2416 54192 -2376
rect 54386 -2416 54406 -2376
rect 54564 -2368 54722 -2358
rect 54564 -2404 54588 -2368
rect 54690 -2404 54722 -2368
rect 54564 -2412 54722 -2404
rect 73858 -2414 73892 -2398
rect 73946 -2170 73980 -2154
rect 73946 -2414 73980 -2398
rect 74076 -2170 74110 -2154
rect 74076 -2414 74110 -2398
rect 74164 -2170 74198 -2154
rect 80446 -2180 80480 -2164
rect 74292 -2278 74374 -2236
rect 74292 -2318 74312 -2278
rect 74350 -2318 74374 -2278
rect 74292 -2344 74374 -2318
rect 80179 -2277 80303 -2242
rect 80179 -2337 80211 -2277
rect 80267 -2337 80303 -2277
rect 80179 -2371 80303 -2337
rect 74164 -2414 74198 -2398
rect 54174 -2432 54406 -2416
rect 80446 -2424 80480 -2408
rect 80534 -2180 80568 -2164
rect 80534 -2424 80568 -2408
rect 80664 -2180 80698 -2164
rect 80664 -2424 80698 -2408
rect 80752 -2180 80786 -2164
rect 99858 -2214 99892 -2198
rect 99946 -1970 99980 -1954
rect 99946 -2214 99980 -2198
rect 100076 -1970 100110 -1954
rect 100076 -2214 100110 -2198
rect 100164 -1970 100198 -1954
rect 106446 -1980 106480 -1964
rect 100342 -2070 100457 -2036
rect 100342 -2122 100370 -2070
rect 100424 -2122 100457 -2070
rect 100342 -2152 100457 -2122
rect 106247 -2097 106346 -2065
rect 106247 -2139 106271 -2097
rect 106313 -2139 106346 -2097
rect 106247 -2161 106346 -2139
rect 100164 -2214 100198 -2198
rect 106446 -2224 106480 -2208
rect 106534 -1980 106568 -1964
rect 106534 -2224 106568 -2208
rect 106664 -1980 106698 -1964
rect 106664 -2224 106698 -2208
rect 106752 -1980 106786 -1964
rect 106752 -2224 106786 -2208
rect 99586 -2266 99818 -2250
rect 99586 -2306 99604 -2266
rect 99798 -2306 99818 -2266
rect 99976 -2258 100134 -2248
rect 99976 -2294 100000 -2258
rect 100102 -2294 100134 -2258
rect 99976 -2302 100134 -2294
rect 106174 -2276 106406 -2260
rect 99586 -2322 99818 -2306
rect 106174 -2316 106192 -2276
rect 106386 -2316 106406 -2276
rect 106564 -2268 106722 -2258
rect 106564 -2304 106588 -2268
rect 106690 -2304 106722 -2268
rect 106564 -2312 106722 -2304
rect 106174 -2332 106406 -2316
rect 80752 -2424 80786 -2408
rect 99858 -2352 99892 -2336
rect 99858 -2428 99892 -2412
rect 99946 -2352 99980 -2336
rect 99946 -2428 99980 -2412
rect 100076 -2352 100110 -2336
rect 100076 -2428 100110 -2412
rect 100164 -2352 100198 -2336
rect 100164 -2428 100198 -2412
rect 106446 -2362 106480 -2346
rect 47858 -2452 47892 -2436
rect 47858 -2528 47892 -2512
rect 47946 -2452 47980 -2436
rect 47946 -2528 47980 -2512
rect 48076 -2452 48110 -2436
rect 48076 -2528 48110 -2512
rect 48164 -2452 48198 -2436
rect 106446 -2438 106480 -2422
rect 106534 -2362 106568 -2346
rect 106534 -2438 106568 -2422
rect 106664 -2362 106698 -2346
rect 106664 -2438 106698 -2422
rect 106752 -2362 106786 -2346
rect 106752 -2438 106786 -2422
rect 48164 -2528 48198 -2512
rect 54446 -2462 54480 -2446
rect 54446 -2538 54480 -2522
rect 54534 -2462 54568 -2446
rect 54534 -2538 54568 -2522
rect 54664 -2462 54698 -2446
rect 54664 -2538 54698 -2522
rect 54752 -2462 54786 -2446
rect 73586 -2466 73818 -2450
rect 73586 -2506 73604 -2466
rect 73798 -2506 73818 -2466
rect 73976 -2458 74134 -2448
rect 73976 -2494 74000 -2458
rect 74102 -2494 74134 -2458
rect 73976 -2502 74134 -2494
rect 80174 -2476 80406 -2460
rect 73586 -2522 73818 -2506
rect 80174 -2516 80192 -2476
rect 80386 -2516 80406 -2476
rect 80564 -2468 80722 -2458
rect 80564 -2504 80588 -2468
rect 80690 -2504 80722 -2468
rect 80564 -2512 80722 -2504
rect 54752 -2538 54786 -2522
rect 80174 -2532 80406 -2516
rect 47258 -2656 47674 -2618
rect 73858 -2552 73892 -2536
rect 73858 -2628 73892 -2612
rect 73946 -2552 73980 -2536
rect 73946 -2628 73980 -2612
rect 74076 -2552 74110 -2536
rect 74076 -2628 74110 -2612
rect 74164 -2552 74198 -2536
rect 74164 -2628 74198 -2612
rect 80446 -2562 80480 -2546
rect 80446 -2638 80480 -2622
rect 80534 -2562 80568 -2546
rect 80534 -2638 80568 -2622
rect 80664 -2562 80698 -2546
rect 80664 -2638 80698 -2622
rect 80752 -2562 80786 -2546
rect 80752 -2638 80786 -2622
<< viali >>
rect 24288 -2216 24324 -2182
rect 30024 -2192 30062 -2156
rect 47332 -2618 47596 -2158
rect 47858 -2298 47892 -2070
rect 47946 -2298 47980 -2070
rect 48076 -2298 48110 -2070
rect 48164 -2298 48198 -2070
rect 48320 -2200 48362 -2164
rect 54304 -2218 54340 -2184
rect 54446 -2308 54480 -2080
rect 54534 -2308 54568 -2080
rect 54664 -2308 54698 -2080
rect 54752 -2308 54786 -2080
rect 48000 -2394 48102 -2358
rect 54192 -2416 54386 -2376
rect 54588 -2404 54690 -2368
rect 73858 -2398 73892 -2170
rect 73946 -2398 73980 -2170
rect 74076 -2398 74110 -2170
rect 74164 -2398 74198 -2170
rect 74312 -2318 74350 -2278
rect 80211 -2337 80267 -2277
rect 80446 -2408 80480 -2180
rect 80534 -2408 80568 -2180
rect 80664 -2408 80698 -2180
rect 80752 -2408 80786 -2180
rect 99858 -2198 99892 -1970
rect 99946 -2198 99980 -1970
rect 100076 -2198 100110 -1970
rect 100164 -2198 100198 -1970
rect 100370 -2122 100424 -2070
rect 106271 -2139 106313 -2097
rect 106446 -2208 106480 -1980
rect 106534 -2208 106568 -1980
rect 106664 -2208 106698 -1980
rect 106752 -2208 106786 -1980
rect 99604 -2306 99798 -2266
rect 100000 -2294 100102 -2258
rect 106192 -2316 106386 -2276
rect 106588 -2304 106690 -2268
rect 99858 -2412 99892 -2352
rect 99946 -2412 99980 -2352
rect 100076 -2412 100110 -2352
rect 100164 -2412 100198 -2352
rect 106446 -2422 106480 -2362
rect 47858 -2512 47892 -2452
rect 47946 -2512 47980 -2452
rect 48076 -2512 48110 -2452
rect 106534 -2422 106568 -2362
rect 106664 -2422 106698 -2362
rect 106752 -2422 106786 -2362
rect 48164 -2512 48198 -2452
rect 54446 -2522 54480 -2462
rect 54534 -2522 54568 -2462
rect 54664 -2522 54698 -2462
rect 54752 -2522 54786 -2462
rect 73604 -2506 73798 -2466
rect 74000 -2494 74102 -2458
rect 80192 -2516 80386 -2476
rect 80588 -2504 80690 -2468
rect 73858 -2612 73892 -2552
rect 73946 -2612 73980 -2552
rect 74076 -2612 74110 -2552
rect 74164 -2612 74198 -2552
rect 80446 -2622 80480 -2562
rect 80534 -2622 80568 -2562
rect 80664 -2622 80698 -2562
rect 80752 -2622 80786 -2562
<< metal1 >>
rect 22480 -1824 30727 -1527
rect 22480 -1997 30738 -1824
rect 22480 -3450 22899 -1997
rect 24288 -2094 24324 -1997
rect 24288 -2158 24326 -2094
rect 30024 -2126 30062 -1997
rect 30302 -2022 30738 -1997
rect 30918 -1888 31702 -1788
rect 29998 -2156 30090 -2126
rect 24264 -2182 24350 -2158
rect 24264 -2216 24288 -2182
rect 24324 -2216 24350 -2182
rect 29998 -2192 30024 -2156
rect 30062 -2192 30090 -2156
rect 29998 -2216 30090 -2192
rect 24264 -2244 24350 -2216
rect 30918 -2366 31002 -1888
rect 24170 -2398 30360 -2370
rect 30808 -2378 31002 -2366
rect 30538 -2406 31002 -2378
rect 23876 -2522 23892 -2518
rect 23858 -2574 23892 -2522
rect 24076 -2574 24110 -2518
rect 30170 -2574 30204 -2526
rect 30388 -2574 30422 -2526
rect 23852 -2584 30438 -2574
rect 30714 -2584 30792 -2574
rect 23852 -2776 30792 -2584
rect 23854 -2942 30792 -2776
rect 30918 -2760 31002 -2406
rect 31590 -2760 31702 -1888
rect 30918 -2842 31702 -2760
rect 46504 -1997 54707 -1750
rect 54922 -1924 55480 -1838
rect 46504 -2003 48111 -1997
rect 22112 -3538 23536 -3450
rect 22112 -3904 22238 -3538
rect 23288 -3904 23536 -3538
rect 22112 -3986 23536 -3904
rect 22695 -3987 22729 -3986
rect 30424 -4302 30792 -2942
rect 46504 -3442 46757 -2003
rect 47858 -2010 48111 -2003
rect 47858 -2058 47892 -2010
rect 48076 -2058 48110 -2010
rect 47852 -2070 47898 -2058
rect 47258 -2158 47674 -2116
rect 47258 -2618 47332 -2158
rect 47596 -2618 47674 -2158
rect 47852 -2298 47858 -2070
rect 47892 -2298 47898 -2070
rect 47852 -2310 47898 -2298
rect 47940 -2070 47986 -2058
rect 47940 -2298 47946 -2070
rect 47980 -2298 47986 -2070
rect 47940 -2310 47986 -2298
rect 48070 -2070 48116 -2058
rect 48070 -2298 48076 -2070
rect 48110 -2298 48116 -2070
rect 48070 -2310 48116 -2298
rect 48158 -2070 48204 -2058
rect 48158 -2298 48164 -2070
rect 48198 -2298 48204 -2070
rect 48320 -2130 48362 -1997
rect 48292 -2164 48394 -2130
rect 54304 -2158 54340 -1997
rect 54446 -2020 54699 -1997
rect 54446 -2068 54480 -2020
rect 54664 -2068 54698 -2020
rect 54440 -2080 54486 -2068
rect 48292 -2200 48320 -2164
rect 48362 -2200 48394 -2164
rect 48292 -2226 48394 -2200
rect 54286 -2184 54358 -2158
rect 54286 -2218 54304 -2184
rect 54340 -2218 54358 -2184
rect 54286 -2246 54358 -2218
rect 48158 -2310 48204 -2298
rect 54440 -2308 54446 -2080
rect 54480 -2308 54486 -2080
rect 47946 -2348 47980 -2310
rect 47946 -2358 48134 -2348
rect 47946 -2394 48000 -2358
rect 48102 -2394 48134 -2358
rect 47946 -2404 48134 -2394
rect 48164 -2370 48198 -2310
rect 54440 -2320 54486 -2308
rect 54528 -2080 54574 -2068
rect 54528 -2308 54534 -2080
rect 54568 -2308 54574 -2080
rect 54528 -2320 54574 -2308
rect 54658 -2080 54704 -2068
rect 54658 -2308 54664 -2080
rect 54698 -2308 54704 -2080
rect 54658 -2320 54704 -2308
rect 54746 -2080 54792 -2068
rect 54746 -2308 54752 -2080
rect 54786 -2308 54792 -2080
rect 54746 -2320 54792 -2308
rect 54534 -2358 54568 -2320
rect 54174 -2368 54406 -2360
rect 54174 -2370 54192 -2368
rect 48164 -2398 54192 -2370
rect 47946 -2440 47980 -2404
rect 48164 -2440 48198 -2398
rect 54174 -2426 54192 -2398
rect 54386 -2426 54406 -2368
rect 54174 -2432 54406 -2426
rect 54534 -2368 54722 -2358
rect 54534 -2404 54588 -2368
rect 54690 -2404 54722 -2368
rect 54534 -2414 54722 -2404
rect 54752 -2366 54786 -2320
rect 54922 -2366 54970 -1924
rect 47852 -2452 47898 -2440
rect 47852 -2512 47858 -2452
rect 47892 -2512 47898 -2452
rect 47852 -2524 47898 -2512
rect 47940 -2452 47986 -2440
rect 47940 -2512 47946 -2452
rect 47980 -2512 47986 -2452
rect 47940 -2524 47986 -2512
rect 48070 -2452 48116 -2440
rect 48070 -2512 48076 -2452
rect 48110 -2512 48116 -2452
rect 48070 -2524 48116 -2512
rect 48158 -2452 48204 -2440
rect 54534 -2450 54568 -2414
rect 54752 -2422 54970 -2366
rect 54752 -2450 54786 -2422
rect 48158 -2512 48164 -2452
rect 48198 -2512 48204 -2452
rect 48158 -2524 48204 -2512
rect 54440 -2462 54486 -2450
rect 54440 -2522 54446 -2462
rect 54480 -2522 54486 -2462
rect 47258 -2656 47674 -2618
rect 47858 -2570 47892 -2524
rect 48076 -2570 48110 -2524
rect 54440 -2534 54486 -2522
rect 54528 -2462 54574 -2450
rect 54528 -2522 54534 -2462
rect 54568 -2522 54574 -2462
rect 54528 -2534 54574 -2522
rect 54658 -2462 54704 -2450
rect 54658 -2522 54664 -2462
rect 54698 -2522 54704 -2462
rect 54658 -2534 54704 -2522
rect 54746 -2462 54792 -2450
rect 54746 -2522 54752 -2462
rect 54786 -2522 54792 -2462
rect 54746 -2534 54792 -2522
rect 54446 -2570 54480 -2534
rect 54664 -2570 54698 -2534
rect 47858 -2573 54846 -2570
rect 47858 -2616 54849 -2573
rect 47858 -2882 54846 -2616
rect 54922 -2764 54970 -2422
rect 55396 -2366 55480 -1924
rect 71998 -2061 80698 -1718
rect 80982 -1930 82012 -1824
rect 71998 -2095 80699 -2061
rect 55396 -2422 55494 -2366
rect 55396 -2764 55480 -2422
rect 54922 -2848 55480 -2764
rect 54534 -3254 54846 -2882
rect 46816 -3442 47111 -3440
rect 46402 -3560 47814 -3442
rect 46402 -3960 46534 -3560
rect 47660 -3960 47814 -3560
rect 46402 -4018 47814 -3960
rect 29948 -4362 31530 -4302
rect 54534 -4322 54849 -3254
rect 71998 -3456 72375 -2095
rect 73858 -2110 74111 -2095
rect 73858 -2158 73892 -2110
rect 74076 -2158 74110 -2110
rect 73096 -2224 73762 -2158
rect 73096 -2776 73186 -2224
rect 73702 -2450 73762 -2224
rect 73852 -2170 73898 -2158
rect 73852 -2398 73858 -2170
rect 73892 -2398 73898 -2170
rect 73852 -2410 73898 -2398
rect 73940 -2170 73986 -2158
rect 73940 -2398 73946 -2170
rect 73980 -2398 73986 -2170
rect 73940 -2410 73986 -2398
rect 74070 -2170 74116 -2158
rect 74070 -2398 74076 -2170
rect 74110 -2398 74116 -2170
rect 74070 -2410 74116 -2398
rect 74158 -2170 74204 -2158
rect 74158 -2398 74164 -2170
rect 74198 -2398 74204 -2170
rect 74312 -2236 74352 -2095
rect 74292 -2278 74374 -2236
rect 80211 -2242 80267 -2095
rect 80446 -2120 80699 -2095
rect 80446 -2168 80480 -2120
rect 80664 -2168 80698 -2120
rect 80440 -2180 80486 -2168
rect 74292 -2318 74312 -2278
rect 74350 -2318 74374 -2278
rect 74292 -2344 74374 -2318
rect 80179 -2277 80303 -2242
rect 80179 -2337 80211 -2277
rect 80267 -2337 80303 -2277
rect 80179 -2371 80303 -2337
rect 74158 -2410 74204 -2398
rect 80440 -2408 80446 -2180
rect 80480 -2408 80486 -2180
rect 73946 -2448 73980 -2410
rect 73702 -2458 73818 -2450
rect 73798 -2516 73818 -2458
rect 73702 -2522 73818 -2516
rect 73946 -2458 74134 -2448
rect 73946 -2494 74000 -2458
rect 74102 -2494 74134 -2458
rect 73946 -2504 74134 -2494
rect 74164 -2470 74198 -2410
rect 80440 -2420 80486 -2408
rect 80528 -2180 80574 -2168
rect 80528 -2408 80534 -2180
rect 80568 -2408 80574 -2180
rect 80528 -2420 80574 -2408
rect 80658 -2180 80704 -2168
rect 80658 -2408 80664 -2180
rect 80698 -2408 80704 -2180
rect 80658 -2420 80704 -2408
rect 80746 -2180 80792 -2168
rect 80746 -2408 80752 -2180
rect 80786 -2408 80792 -2180
rect 80746 -2420 80792 -2408
rect 80534 -2458 80568 -2420
rect 80174 -2468 80406 -2460
rect 80174 -2470 80192 -2468
rect 74164 -2498 80192 -2470
rect 73702 -2776 73762 -2522
rect 73946 -2540 73980 -2504
rect 74164 -2540 74198 -2498
rect 80174 -2526 80192 -2498
rect 80386 -2526 80406 -2468
rect 80174 -2532 80406 -2526
rect 80534 -2468 80722 -2458
rect 80534 -2504 80588 -2468
rect 80690 -2504 80722 -2468
rect 80534 -2514 80722 -2504
rect 80752 -2466 80786 -2420
rect 80982 -2466 81084 -1930
rect 73852 -2552 73898 -2540
rect 73852 -2612 73858 -2552
rect 73892 -2612 73898 -2552
rect 73852 -2624 73898 -2612
rect 73940 -2552 73986 -2540
rect 73940 -2612 73946 -2552
rect 73980 -2612 73986 -2552
rect 73940 -2624 73986 -2612
rect 74070 -2552 74116 -2540
rect 74070 -2612 74076 -2552
rect 74110 -2612 74116 -2552
rect 74070 -2624 74116 -2612
rect 74158 -2552 74204 -2540
rect 80534 -2550 80568 -2514
rect 80752 -2522 81084 -2466
rect 80752 -2550 80786 -2522
rect 74158 -2612 74164 -2552
rect 74198 -2612 74204 -2552
rect 74158 -2624 74204 -2612
rect 80440 -2562 80486 -2550
rect 80440 -2622 80446 -2562
rect 80480 -2622 80486 -2562
rect 73858 -2689 73892 -2624
rect 74076 -2689 74110 -2624
rect 80440 -2634 80486 -2622
rect 80528 -2562 80574 -2550
rect 80528 -2622 80534 -2562
rect 80568 -2622 80574 -2562
rect 80528 -2634 80574 -2622
rect 80658 -2562 80704 -2550
rect 80658 -2622 80664 -2562
rect 80698 -2622 80704 -2562
rect 80658 -2634 80704 -2622
rect 80746 -2562 80792 -2550
rect 80746 -2622 80752 -2562
rect 80786 -2622 80792 -2562
rect 80746 -2634 80792 -2622
rect 80446 -2689 80480 -2634
rect 80664 -2689 80698 -2634
rect 73858 -2692 80867 -2689
rect 73096 -2846 73762 -2776
rect 73850 -2976 80867 -2692
rect 80982 -2768 81084 -2522
rect 81850 -2768 82012 -1930
rect 80982 -2846 82012 -2768
rect 97086 -1898 106786 -1538
rect 72448 -3456 72804 -3436
rect 71904 -3538 73800 -3456
rect 71904 -3896 72176 -3538
rect 73580 -3896 73800 -3538
rect 71904 -3990 73800 -3896
rect 80580 -4294 80867 -2976
rect 97086 -3456 97446 -1898
rect 99858 -1910 100111 -1898
rect 99858 -1958 99892 -1910
rect 100076 -1958 100110 -1910
rect 99852 -1970 99898 -1958
rect 99852 -2198 99858 -1970
rect 99892 -2198 99898 -1970
rect 99852 -2210 99898 -2198
rect 99940 -1970 99986 -1958
rect 99940 -2198 99946 -1970
rect 99980 -2198 99986 -1970
rect 99940 -2210 99986 -2198
rect 100070 -1970 100116 -1958
rect 100070 -2198 100076 -1970
rect 100110 -2198 100116 -1970
rect 100070 -2210 100116 -2198
rect 100158 -1970 100204 -1958
rect 100158 -2198 100164 -1970
rect 100198 -2198 100204 -1970
rect 100370 -2036 100424 -1898
rect 100342 -2070 100457 -2036
rect 106270 -2065 106315 -1898
rect 106446 -1920 106699 -1898
rect 106446 -1968 106480 -1920
rect 106664 -1968 106698 -1920
rect 107068 -1952 107998 -1768
rect 106440 -1980 106486 -1968
rect 100342 -2122 100370 -2070
rect 100424 -2122 100457 -2070
rect 100342 -2152 100457 -2122
rect 106247 -2097 106346 -2065
rect 106247 -2139 106271 -2097
rect 106313 -2139 106346 -2097
rect 106247 -2161 106346 -2139
rect 100158 -2210 100204 -2198
rect 106440 -2208 106446 -1980
rect 106480 -2208 106486 -1980
rect 99946 -2248 99980 -2210
rect 99586 -2258 99818 -2250
rect 99586 -2316 99604 -2258
rect 99798 -2316 99818 -2258
rect 99586 -2322 99818 -2316
rect 99946 -2258 100134 -2248
rect 99946 -2294 100000 -2258
rect 100102 -2294 100134 -2258
rect 99946 -2304 100134 -2294
rect 100164 -2270 100198 -2210
rect 106440 -2220 106486 -2208
rect 106528 -1980 106574 -1968
rect 106528 -2208 106534 -1980
rect 106568 -2208 106574 -1980
rect 106528 -2220 106574 -2208
rect 106658 -1980 106704 -1968
rect 106658 -2208 106664 -1980
rect 106698 -2208 106704 -1980
rect 106658 -2220 106704 -2208
rect 106746 -1980 106792 -1968
rect 106746 -2208 106752 -1980
rect 106786 -2208 106792 -1980
rect 106746 -2220 106792 -2208
rect 106534 -2258 106568 -2220
rect 106174 -2268 106406 -2260
rect 106174 -2270 106192 -2268
rect 100164 -2298 106192 -2270
rect 99946 -2340 99980 -2304
rect 100164 -2340 100198 -2298
rect 106174 -2326 106192 -2298
rect 106386 -2326 106406 -2268
rect 106174 -2332 106406 -2326
rect 106534 -2268 106722 -2258
rect 106534 -2304 106588 -2268
rect 106690 -2304 106722 -2268
rect 106534 -2314 106722 -2304
rect 106752 -2266 106786 -2220
rect 107068 -2266 107200 -1952
rect 99852 -2352 99898 -2340
rect 99852 -2412 99858 -2352
rect 99892 -2412 99898 -2352
rect 99852 -2424 99898 -2412
rect 99940 -2352 99986 -2340
rect 99940 -2412 99946 -2352
rect 99980 -2412 99986 -2352
rect 99940 -2424 99986 -2412
rect 100070 -2352 100116 -2340
rect 100070 -2412 100076 -2352
rect 100110 -2412 100116 -2352
rect 100070 -2424 100116 -2412
rect 100158 -2352 100204 -2340
rect 106534 -2350 106568 -2314
rect 106752 -2322 107200 -2266
rect 106752 -2350 106786 -2322
rect 100158 -2412 100164 -2352
rect 100198 -2412 100204 -2352
rect 100158 -2424 100204 -2412
rect 106440 -2362 106486 -2350
rect 106440 -2422 106446 -2362
rect 106480 -2422 106486 -2362
rect 99858 -2513 99892 -2424
rect 100076 -2513 100110 -2424
rect 106440 -2434 106486 -2422
rect 106528 -2362 106574 -2350
rect 106528 -2422 106534 -2362
rect 106568 -2422 106574 -2362
rect 106528 -2434 106574 -2422
rect 106658 -2362 106704 -2350
rect 106658 -2422 106664 -2362
rect 106698 -2422 106704 -2362
rect 106658 -2434 106704 -2422
rect 106746 -2362 106792 -2350
rect 106746 -2422 106752 -2362
rect 106786 -2422 106792 -2362
rect 106746 -2434 106792 -2422
rect 106446 -2513 106480 -2434
rect 106664 -2513 106698 -2434
rect 99858 -2524 106841 -2513
rect 99842 -2640 106841 -2524
rect 99850 -2836 106841 -2640
rect 96740 -3524 98336 -3456
rect 96740 -3922 96888 -3524
rect 98194 -3922 98336 -3524
rect 96740 -4006 98336 -3922
rect 97086 -4022 97446 -4006
rect 29948 -4824 30068 -4362
rect 31382 -4824 31530 -4362
rect 29948 -4888 31530 -4824
rect 53726 -4426 55902 -4322
rect 53726 -4796 53860 -4426
rect 55650 -4796 55902 -4426
rect 53726 -4878 55902 -4796
rect 80010 -4364 81428 -4294
rect 80010 -4830 80140 -4364
rect 81300 -4830 81428 -4364
rect 54815 -4885 54849 -4878
rect 30561 -4897 30763 -4888
rect 80010 -4890 81428 -4830
rect 106094 -4296 106266 -4292
rect 106518 -4296 106841 -2836
rect 107068 -2742 107200 -2322
rect 107808 -2742 107998 -1952
rect 107068 -2850 107998 -2742
rect 106094 -4390 107330 -4296
rect 106094 -4838 106210 -4390
rect 107214 -4838 107330 -4390
rect 80694 -4907 80841 -4890
rect 106094 -4894 107330 -4838
<< via1 >>
rect 31002 -2760 31590 -1888
rect 22238 -3904 23288 -3538
rect 47332 -2618 47596 -2158
rect 54192 -2376 54386 -2368
rect 54192 -2416 54386 -2376
rect 54192 -2426 54386 -2416
rect 54970 -2764 55396 -1924
rect 46534 -3960 47660 -3560
rect 73186 -2458 73702 -2224
rect 73186 -2466 73798 -2458
rect 73186 -2506 73604 -2466
rect 73604 -2506 73798 -2466
rect 73186 -2516 73798 -2506
rect 73186 -2776 73702 -2516
rect 80192 -2476 80386 -2468
rect 80192 -2516 80386 -2476
rect 80192 -2526 80386 -2516
rect 81084 -2768 81850 -1930
rect 72176 -3896 73580 -3538
rect 99604 -2266 99798 -2258
rect 99604 -2306 99798 -2266
rect 99604 -2316 99798 -2306
rect 106192 -2276 106386 -2268
rect 106192 -2316 106386 -2276
rect 106192 -2326 106386 -2316
rect 96888 -3922 98194 -3524
rect 30068 -4824 31382 -4362
rect 53860 -4796 55650 -4426
rect 80140 -4830 81300 -4364
rect 107200 -2742 107808 -1952
rect 106210 -4838 107214 -4390
<< metal2 >>
rect 50889 25140 51036 25224
rect 102471 25156 102614 25240
rect 50952 24592 51036 25140
rect 102530 24616 102614 25156
rect 23952 23380 27286 23440
rect 49356 23402 52704 23468
rect 74898 23394 78854 23458
rect 100930 23420 104262 23480
rect 23934 21288 27268 21348
rect 49318 21292 52666 21358
rect 74894 21296 78850 21360
rect 100900 21316 104232 21376
rect 23902 19194 27236 19254
rect 49336 19196 52684 19262
rect 74872 19204 78828 19268
rect 100930 19214 104262 19274
rect 23960 17096 27294 17156
rect 49400 17098 52748 17164
rect 74908 17112 78864 17176
rect 100980 17128 104312 17188
rect 23916 15004 27250 15064
rect 49450 15010 52798 15076
rect 74882 15022 78838 15086
rect 101012 15034 104344 15094
rect 23844 12910 27280 12970
rect 49388 12918 52736 12984
rect 74830 12926 78854 12994
rect 100972 12938 104328 13002
rect 23820 10816 27294 10872
rect 49416 10834 52702 10874
rect 74828 10838 78852 10906
rect 100986 10848 104342 10912
rect 23816 8716 27290 8772
rect 49562 8730 52622 8792
rect 74808 8730 78878 8800
rect 100992 8738 104348 8802
rect 25458 7020 25542 7594
rect 77072 7042 77156 7608
rect 25362 6936 25542 7020
rect 76364 6958 77156 7042
rect 30918 -1888 31702 -1788
rect 23136 -2238 23664 -2150
rect 23136 -2796 23210 -2238
rect 23570 -2796 23664 -2238
rect 23136 -2846 23664 -2796
rect 30918 -2760 31002 -1888
rect 31590 -2760 31702 -1888
rect 54922 -1924 55480 -1838
rect 47258 -2158 47674 -2116
rect 47258 -2618 47332 -2158
rect 47596 -2618 47674 -2158
rect 54174 -2368 54406 -2360
rect 54174 -2426 54192 -2368
rect 54386 -2426 54406 -2368
rect 54174 -2432 54406 -2426
rect 47258 -2656 47674 -2618
rect 30918 -2842 31702 -2760
rect 54922 -2764 54970 -1924
rect 55396 -2764 55480 -1924
rect 80982 -1930 82012 -1824
rect 54922 -2848 55480 -2764
rect 73096 -2224 73772 -2158
rect 73096 -2776 73186 -2224
rect 73702 -2442 73772 -2224
rect 73702 -2450 73816 -2442
rect 73702 -2458 73818 -2450
rect 73798 -2516 73818 -2458
rect 73702 -2522 73818 -2516
rect 80174 -2468 80406 -2460
rect 73702 -2530 73816 -2522
rect 80174 -2526 80192 -2468
rect 80386 -2526 80406 -2468
rect 73702 -2776 73772 -2530
rect 80174 -2532 80406 -2526
rect 73096 -2846 73772 -2776
rect 80982 -2768 81084 -1930
rect 81850 -2768 82012 -1930
rect 107068 -1952 107998 -1768
rect 80982 -2846 82012 -2768
rect 99190 -2142 99764 -2058
rect 99190 -2776 99256 -2142
rect 99696 -2242 99764 -2142
rect 99696 -2250 99816 -2242
rect 99696 -2258 99818 -2250
rect 99798 -2316 99818 -2258
rect 99696 -2322 99818 -2316
rect 106174 -2268 106406 -2260
rect 99696 -2330 99816 -2322
rect 106174 -2326 106192 -2268
rect 106386 -2326 106406 -2268
rect 99696 -2776 99764 -2330
rect 106174 -2332 106406 -2326
rect 99190 -2824 99764 -2776
rect 107068 -2742 107200 -1952
rect 107808 -2742 107998 -1952
rect 107068 -2850 107998 -2742
rect 22112 -3538 23536 -3450
rect 22112 -3904 22238 -3538
rect 23288 -3904 23536 -3538
rect 22112 -3986 23536 -3904
rect 46402 -3560 47814 -3442
rect 46402 -3960 46534 -3560
rect 47660 -3960 47814 -3560
rect 46402 -4018 47814 -3960
rect 71904 -3538 73800 -3456
rect 71904 -3896 72176 -3538
rect 73580 -3896 73800 -3538
rect 71904 -3990 73800 -3896
rect 96740 -3524 98336 -3456
rect 96740 -3922 96888 -3524
rect 98194 -3922 98336 -3524
rect 96740 -4006 98336 -3922
rect 29948 -4362 31530 -4302
rect 29948 -4824 30068 -4362
rect 31382 -4824 31530 -4362
rect 29948 -4888 31530 -4824
rect 53726 -4426 55902 -4322
rect 53726 -4796 53860 -4426
rect 55650 -4796 55902 -4426
rect 53726 -4878 55902 -4796
rect 80010 -4364 81428 -4294
rect 80010 -4830 80140 -4364
rect 81300 -4830 81428 -4364
rect 80010 -4890 81428 -4830
rect 106094 -4296 106266 -4292
rect 106094 -4390 107330 -4296
rect 106094 -4838 106210 -4390
rect 107214 -4838 107330 -4390
rect 106094 -4894 107330 -4838
<< via2 >>
rect 23210 -2796 23570 -2238
rect 31002 -2760 31590 -1888
rect 47332 -2618 47596 -2158
rect 54970 -2764 55396 -1924
rect 73186 -2776 73702 -2224
rect 81084 -2768 81850 -1930
rect 99256 -2258 99696 -2142
rect 99256 -2316 99604 -2258
rect 99604 -2316 99696 -2258
rect 99256 -2776 99696 -2316
rect 107200 -2742 107808 -1952
rect 22238 -3904 23288 -3538
rect 46534 -3960 47660 -3560
rect 72176 -3896 73580 -3538
rect 96888 -3922 98194 -3524
rect 30068 -4824 31382 -4362
rect 53860 -4796 55650 -4426
rect 80140 -4830 81300 -4364
rect 106210 -4838 107214 -4390
<< metal3 >>
rect 12789 -1800 12923 134
rect 38498 -1800 38570 -1048
rect 63771 -1800 63905 156
rect 90070 -1800 90142 -1026
rect 115359 -1800 115493 231
rect -1718 -2238 23667 -1800
rect -1718 -2796 23210 -2238
rect 23570 -2796 23667 -2238
rect -1718 -2858 23667 -2796
rect 30907 -1888 47685 -1800
rect 30907 -2760 31002 -1888
rect 31590 -2158 47685 -1888
rect 31590 -2618 47332 -2158
rect 47596 -2618 47685 -2158
rect 31590 -2760 47685 -2618
rect 30907 -2858 47685 -2760
rect 54901 -1924 73833 -1800
rect 54901 -2764 54970 -1924
rect 55396 -2224 73833 -1924
rect 55396 -2764 73186 -2224
rect 54901 -2776 73186 -2764
rect 73702 -2776 73833 -2224
rect 54901 -2858 73833 -2776
rect 80965 -1930 99801 -1800
rect 80965 -2768 81084 -1930
rect 81850 -2142 99801 -1930
rect 81850 -2768 99256 -2142
rect 80965 -2776 99256 -2768
rect 99696 -2776 99801 -2142
rect 80965 -2858 99801 -2776
rect 106853 -1952 115780 -1800
rect 106853 -2742 107200 -1952
rect 107808 -2742 115780 -1952
rect 106853 -2858 115780 -2742
rect 22112 -3538 23536 -3450
rect 22112 -3904 22238 -3538
rect 23288 -3904 23536 -3538
rect 22112 -3986 23536 -3904
rect 46402 -3560 47814 -3442
rect 46402 -3960 46534 -3560
rect 47660 -3960 47814 -3560
rect 46402 -4018 47814 -3960
rect 71904 -3538 73800 -3456
rect 71904 -3896 72176 -3538
rect 73580 -3896 73800 -3538
rect 71904 -3990 73800 -3896
rect 96740 -3524 98336 -3456
rect 96740 -3922 96888 -3524
rect 98194 -3922 98336 -3524
rect 96740 -4006 98336 -3922
rect 29948 -4362 31530 -4302
rect 29948 -4824 30068 -4362
rect 31382 -4824 31530 -4362
rect 29948 -4888 31530 -4824
rect 53726 -4426 55902 -4322
rect 53726 -4796 53860 -4426
rect 55650 -4796 55902 -4426
rect 53726 -4878 55902 -4796
rect 80010 -4364 81428 -4294
rect 80010 -4830 80140 -4364
rect 81300 -4830 81428 -4364
rect 80010 -4890 81428 -4830
rect 106094 -4296 106266 -4292
rect 106094 -4390 107330 -4296
rect 106094 -4838 106210 -4390
rect 107214 -4838 107330 -4390
rect 106094 -4894 107330 -4838
<< via3 >>
rect 22238 -3904 23288 -3538
rect 46534 -3960 47660 -3560
rect 72176 -3896 73580 -3538
rect 96888 -3922 98194 -3524
rect 30068 -4824 31382 -4362
rect 53860 -4796 55650 -4426
rect 80140 -4830 81300 -4364
rect 106210 -4838 107214 -4390
<< metal4 >>
rect 980 -3440 1548 2756
rect 43966 -3440 44550 3340
rect 59884 -3440 60452 2554
rect 95684 -3440 96268 3806
rect 112564 -3440 113132 2522
rect 980 -3524 113132 -3440
rect 980 -3538 96888 -3524
rect 980 -3904 22238 -3538
rect 23288 -3560 72176 -3538
rect 23288 -3904 46534 -3560
rect 980 -3960 46534 -3904
rect 47660 -3896 72176 -3560
rect 73580 -3896 96888 -3538
rect 47660 -3922 96888 -3896
rect 98194 -3922 113132 -3524
rect 47660 -3960 113132 -3922
rect 980 -4008 113132 -3960
rect 43966 -4074 44550 -4008
rect 46402 -4018 47814 -4008
rect 29948 -4362 31530 -4302
rect 29948 -4824 30068 -4362
rect 31382 -4824 31530 -4362
rect 29948 -4888 31530 -4824
rect 53726 -4426 55902 -4322
rect 53726 -4796 53860 -4426
rect 55650 -4796 55902 -4426
rect 53726 -4878 55902 -4796
rect 80010 -4364 81428 -4294
rect 80010 -4830 80140 -4364
rect 81300 -4830 81428 -4364
rect 80010 -4890 81428 -4830
rect 106094 -4296 106266 -4292
rect 106094 -4390 107330 -4296
rect 106094 -4838 106210 -4390
rect 107214 -4838 107330 -4390
rect 106094 -4894 107330 -4838
<< via4 >>
rect 30068 -4824 31382 -4362
rect 53860 -4796 55650 -4426
rect 80140 -4830 81300 -4364
rect 106210 -4838 107214 -4390
<< metal5 >>
rect 281 -4294 885 8386
rect 17957 -4294 18547 2893
rect 34625 -4294 35215 3705
rect 69705 -4294 70295 2915
rect 86083 -4294 86673 3721
rect 127376 -4294 127966 3435
rect 281 -4296 106266 -4294
rect 107746 -4296 128160 -4294
rect 281 -4362 128160 -4296
rect 281 -4824 30068 -4362
rect 31382 -4364 128160 -4362
rect 31382 -4426 80140 -4364
rect 31382 -4796 53860 -4426
rect 55650 -4796 80140 -4426
rect 31382 -4824 80140 -4796
rect 281 -4830 80140 -4824
rect 81300 -4390 128160 -4364
rect 81300 -4830 106210 -4390
rect 281 -4838 106210 -4830
rect 107214 -4838 128160 -4390
rect 281 -4898 128160 -4838
use buffer_digital  buffer_digital_0 ~/Desktop/charge_pumps2/layout_files
timestamp 1698753667
transform 1 0 23860 0 1 -2552
box -274 0 415 576
use buffer_digital  buffer_digital_1
timestamp 1698753667
transform 1 0 30172 0 1 -2560
box -274 0 415 576
use charge_pump1  charge_pump1_0
timestamp 1698753667
transform 1 0 313 0 1 7588
box -313 -7588 25321 19132
use charge_pump1  charge_pump1_1
timestamp 1698753667
transform 1 0 51295 0 1 7610
box -313 -7588 25321 19132
use charge_pump1  charge_pump1_2
timestamp 1698753667
transform 1 0 102883 0 1 7632
box -313 -7588 25321 19132
use charge_pump1_reverse  charge_pump1_reverse_0
timestamp 1698753667
transform 1 0 25809 0 -1 24570
box -313 -3396 25321 25896
use charge_pump1_reverse  charge_pump1_reverse_1
timestamp 1698753667
transform 1 0 77391 0 -1 24582
box -313 -3396 25321 25896
<< end >>
