magic
tech sky130A
magscale 1 2
timestamp 1698869963
<< nwell >>
rect 30476 -606 37144 -32
rect 38102 -732 38770 -490
rect 41350 -746 50272 -46
rect 37634 -1454 39158 -1118
<< nsubdiff >>
rect 38274 -560 38508 -534
rect 38274 -658 38310 -560
rect 38462 -658 38508 -560
rect 38274 -682 38508 -658
<< nsubdiffcont >>
rect 38310 -658 38462 -560
<< locali >>
rect 38274 -560 38508 -534
rect 38274 -658 38310 -560
rect 38462 -658 38508 -560
rect 38274 -682 38508 -658
<< viali >>
rect 38310 -658 38462 -560
<< metal1 >>
rect 28380 -1218 28820 8648
rect 29004 6800 29424 6812
rect 29004 6752 29446 6800
rect 29004 6096 29078 6752
rect 29394 6096 29446 6752
rect 29004 6052 29446 6096
rect 29012 3660 29446 6052
rect 29012 3236 29474 3660
rect 29022 76 29474 3236
rect 50136 76 50510 6760
rect 29022 -222 50510 76
rect 29022 -328 37806 -222
rect 37742 -448 37806 -328
rect 39112 -328 50510 -222
rect 39112 -448 39200 -328
rect 50136 -346 50510 -328
rect 29590 -1218 37096 -462
rect 37742 -478 39200 -448
rect 38274 -560 38512 -478
rect 38274 -658 38310 -560
rect 38462 -658 38512 -560
rect 38274 -682 38512 -658
rect 39468 -590 39790 -558
rect 39468 -840 39498 -590
rect 38117 -883 38606 -850
rect 39175 -873 39498 -840
rect 39468 -890 39498 -873
rect 39746 -890 39790 -590
rect 39468 -940 39790 -890
rect 37742 -1118 37776 -996
rect 37960 -1118 37994 -996
rect 38800 -1118 38834 -986
rect 39018 -1118 39052 -985
rect 37634 -1168 39158 -1118
rect 37634 -1218 37754 -1168
rect 28380 -1416 37754 -1218
rect 39040 -1218 39158 -1168
rect 40490 -1218 49412 -554
rect 50708 -1218 51110 7884
rect 39040 -1416 51130 -1218
rect 28380 -1688 51130 -1416
<< via1 >>
rect 29078 6096 29394 6752
rect 37806 -448 39112 -222
rect 39498 -890 39746 -590
rect 37754 -1416 39040 -1168
<< metal2 >>
rect 29004 6752 29424 6812
rect 29004 6096 29078 6752
rect 29394 6096 29424 6752
rect 29004 6052 29424 6096
rect 37746 -222 39196 -186
rect 37746 -448 37806 -222
rect 39112 -448 39196 -222
rect 37746 -468 39196 -448
rect 37248 -598 37648 -568
rect 37248 -900 37296 -598
rect 37558 -900 37648 -598
rect 37248 -936 37648 -900
rect 39468 -590 39790 -558
rect 39468 -890 39498 -590
rect 39746 -890 39790 -590
rect 39468 -940 39790 -890
rect 37634 -1168 39158 -1118
rect 37634 -1416 37754 -1168
rect 39040 -1416 39158 -1168
rect 37634 -1454 39158 -1416
<< via2 >>
rect 29078 6096 29394 6752
rect 37806 -448 39112 -222
rect 37296 -900 37558 -598
rect 39498 -890 39746 -590
rect 37754 -1416 39040 -1168
<< metal3 >>
rect 29004 6752 29424 6812
rect 29004 6096 29078 6752
rect 29394 6096 29424 6752
rect 29004 6052 29424 6096
rect 37742 -222 39200 -188
rect 37742 -448 37806 -222
rect 39112 -448 39200 -222
rect 37742 -478 39200 -448
rect 39964 -554 40036 770
rect 28014 -598 37654 -556
rect 28014 -900 37296 -598
rect 37558 -900 37654 -598
rect 28014 -948 37654 -900
rect 39456 -590 50472 -554
rect 39456 -890 39498 -590
rect 39746 -890 50472 -590
rect 39456 -946 50472 -890
rect 37632 -1168 39152 -1118
rect 37632 -1416 37754 -1168
rect 39040 -1416 39152 -1168
rect 37632 -1454 39152 -1416
<< via3 >>
rect 29078 6096 29394 6752
rect 37806 -448 39112 -222
rect 37754 -1416 39040 -1168
<< metal4 >>
rect 28903 6752 29601 10459
rect 28903 6096 29078 6752
rect 29394 6096 29601 6752
rect 28903 225 29601 6096
rect 50708 5073 51110 7884
rect 50078 225 51110 5073
rect 28014 -222 51110 225
rect 28014 -448 37806 -222
rect 39112 -448 51110 -222
rect 28014 -473 51110 -448
rect 37634 -1168 39158 -1118
rect 37634 -1416 37754 -1168
rect 39040 -1416 39158 -1168
rect 37634 -1454 39158 -1416
rect 50708 -1668 51110 -473
<< via4 >>
rect 37754 -1416 39040 -1168
<< metal5 >>
rect 28272 -1088 28930 4791
rect 50606 -1088 51264 10087
rect 28014 -1168 51269 -1088
rect 28014 -1416 37754 -1168
rect 39040 -1416 51269 -1168
rect 28014 -1767 51269 -1416
rect 50606 -1775 51264 -1767
use buffer_digital  buffer_digital_2 ~/Desktop/charge_pumps2/layout_files
timestamp 1698771642
transform 1 0 37744 0 1 -1030
box -274 0 415 576
use buffer_digital  buffer_digital_3
timestamp 1698771642
transform 1 0 38802 0 1 -1020
box -274 0 415 576
use charge_pump_reverse  charge_pump_reverse_0
timestamp 1698849032
transform 1 0 27508 0 -1 26452
box 498 -3206 23756 25968
use nmos_decap_10  nmos_decap_10_0
timestamp 1698837560
transform 0 1 28776 -1 0 1188
box -10 -42 1060 416
use nmos_decap_10  nmos_decap_10_1
timestamp 1698837560
transform 0 1 28776 -1 0 2148
box -10 -42 1060 416
use nmos_decap_10  nmos_decap_10_2
timestamp 1698837560
transform 0 1 28776 -1 0 3108
box -10 -42 1060 416
use nmos_decap_10  nmos_decap_10_3
timestamp 1698837560
transform 0 1 28776 -1 0 4068
box -10 -42 1060 416
use nmos_decap_10  nmos_decap_10_4
timestamp 1698837560
transform 0 1 28776 -1 0 5028
box -10 -42 1060 416
use nmos_decap_10  nmos_decap_10_5
timestamp 1698837560
transform 0 1 28776 -1 0 5988
box -10 -42 1060 416
use nmos_decap_10  nmos_decap_10_6
timestamp 1698837560
transform 0 -1 50756 -1 0 1266
box -10 -42 1060 416
use nmos_decap_10  nmos_decap_10_7
timestamp 1698837560
transform 0 -1 50756 -1 0 2226
box -10 -42 1060 416
use nmos_decap_10  nmos_decap_10_8
timestamp 1698837560
transform 0 -1 50756 -1 0 3186
box -10 -42 1060 416
use nmos_decap_10  nmos_decap_10_9
timestamp 1698837560
transform 0 -1 50756 -1 0 4146
box -10 -42 1060 416
use pmos_decap_10  pmos_decap_10_0
timestamp 1698841269
transform 1 0 29506 0 -1 -142
box 0 -108 1098 464
use pmos_decap_10  pmos_decap_10_1
timestamp 1698841269
transform 1 0 30578 0 -1 -134
box 0 -108 1098 464
use pmos_decap_10  pmos_decap_10_2
timestamp 1698841269
transform 1 0 31652 0 -1 -138
box 0 -108 1098 464
use pmos_decap_10  pmos_decap_10_3
timestamp 1698841269
transform 1 0 32724 0 -1 -136
box 0 -108 1098 464
use pmos_decap_10  pmos_decap_10_4
timestamp 1698841269
transform 1 0 33798 0 -1 -140
box 0 -108 1098 464
use pmos_decap_10  pmos_decap_10_5
timestamp 1698841269
transform 1 0 34872 0 -1 -140
box 0 -108 1098 464
use pmos_decap_10  pmos_decap_10_6
timestamp 1698841269
transform 1 0 35944 0 -1 -138
box 0 -108 1098 464
use pmos_decap_10  pmos_decap_10_7
timestamp 1698841269
transform 1 0 40458 0 -1 -146
box 0 -108 1098 464
use pmos_decap_10  pmos_decap_10_8
timestamp 1698841269
transform 1 0 41530 0 -1 -146
box 0 -108 1098 464
use pmos_decap_10  pmos_decap_10_9
timestamp 1698841269
transform 1 0 42602 0 -1 -142
box 0 -108 1098 464
use pmos_decap_10  pmos_decap_10_10
timestamp 1698841269
transform 1 0 43674 0 -1 -146
box 0 -108 1098 464
use pmos_decap_10  pmos_decap_10_11
timestamp 1698841269
transform 1 0 44748 0 -1 -142
box 0 -108 1098 464
use pmos_decap_10  pmos_decap_10_12
timestamp 1698841269
transform 1 0 45820 0 -1 -146
box 0 -108 1098 464
use pmos_decap_10  pmos_decap_10_13
timestamp 1698841269
transform 1 0 46894 0 -1 -146
box 0 -108 1098 464
use pmos_decap_10  pmos_decap_10_14
timestamp 1698841269
transform 1 0 47966 0 -1 -142
box 0 -108 1098 464
use pmos_decap_10  pmos_decap_10_15
timestamp 1698841269
transform 1 0 49038 0 -1 -142
box 0 -108 1098 464
<< end >>
