* SPICE3 file created from reconfigurable_CP.ext - technology: sky130A

.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
X0 VPWR VGND VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0.452 ps=4.52 w=0.87 l=0.59
X1 VGND VPWR VGND VNB sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0.286 ps=3.24 w=0.55 l=0.59
.ends

.subckt sky130_fd_sc_hd__a21oi_1 A1 A2 B1 VGND VNB VPB VPWR Y
X0 a_199_47# A1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.0959 pd=0.945 as=0.091 ps=0.93 w=0.65 l=0.15
X1 a_113_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.147 ps=1.29 w=1 l=0.15
X2 Y B1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.172 ps=1.83 w=0.65 l=0.15
X3 VPWR A1 a_113_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.147 pd=1.29 as=0.14 ps=1.28 w=1 l=0.15
X4 a_113_297# B1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X5 VGND A2 a_199_47# VNB sky130_fd_pr__nfet_01v8 ad=0.172 pd=1.83 as=0.0959 ps=0.945 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__o31a_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
X0 a_103_199# B1 a_253_47# VNB sky130_fd_pr__nfet_01v8 ad=0.201 pd=1.92 as=0.107 ps=0.98 w=0.65 l=0.15
X1 VPWR a_103_199# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=1.39 as=0.36 ps=2.72 w=1 l=0.15
X2 a_337_297# A2 a_253_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.135 ps=1.27 w=1 l=0.15
X3 a_103_199# A3 a_337_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.213 pd=1.42 as=0.165 ps=1.33 w=1 l=0.15
X4 a_253_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.195 ps=1.39 w=1 l=0.15
X5 VPWR B1 a_103_199# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.345 pd=2.69 as=0.213 ps=1.42 w=1 l=0.15
X6 VGND a_103_199# X VNB sky130_fd_pr__nfet_01v8 ad=0.127 pd=1.04 as=0.234 ps=2.02 w=0.65 l=0.15
X7 a_253_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.127 ps=1.04 w=0.65 l=0.15
X8 a_253_47# A3 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.107 ps=0.98 w=0.65 l=0.15
X9 VGND A2 a_253_47# VNB sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.0878 ps=0.92 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
X0 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X1 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.149 ps=1.33 w=1 l=0.15
X2 VPWR A a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.33 as=0.166 ps=1.8 w=0.64 l=0.15
X3 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X4 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.172 pd=1.83 as=0.0878 ps=0.92 w=0.65 l=0.15
X5 VGND A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__or3_1 A B C VGND VNB VPB VPWR X
X0 X a_29_53# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.148 ps=1.34 w=1 l=0.15
X1 a_111_297# C a_29_53# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.109 ps=1.36 w=0.42 l=0.15
X2 X a_29_53# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.102 ps=0.99 w=0.65 l=0.15
X3 a_183_297# B a_111_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X4 VPWR A a_183_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.148 pd=1.34 as=0.0693 ps=0.75 w=0.42 l=0.15
X5 a_29_53# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X6 VGND C a_29_53# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X7 VGND A a_29_53# VNB sky130_fd_pr__nfet_01v8 ad=0.102 pd=0.99 as=0.0567 ps=0.69 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__clkbuf_4 A VGND VNB VPB VPWR X
X0 VPWR A a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.265 ps=2.53 w=1 l=0.15
X1 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0588 ps=0.7 w=0.42 l=0.15
X2 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X5 VGND A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0703 pd=0.755 as=0.111 ps=1.37 w=0.42 l=0.15
X6 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.14 ps=1.28 w=1 l=0.15
X7 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0703 ps=0.755 w=0.42 l=0.15
X8 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.165 ps=1.33 w=1 l=0.15
X9 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
.ends

.subckt sky130_fd_sc_hd__o21a_1 A1 A2 B1 VGND VNB VPB VPWR X
X0 VPWR A1 a_382_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.153 ps=1.3 w=1 l=0.15
X1 a_297_47# B1 a_79_21# VNB sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.96 as=0.169 ps=1.82 w=0.65 l=0.15
X2 a_297_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X3 VGND A2 a_297_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.101 ps=0.96 w=0.65 l=0.15
X4 VPWR a_79_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.327 pd=1.65 as=0.28 ps=2.56 w=1 l=0.15
X5 a_79_21# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=1.39 as=0.327 ps=1.65 w=1 l=0.15
X6 a_382_297# A2 a_79_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.153 pd=1.3 as=0.195 ps=1.39 w=1 l=0.15
X7 VGND a_79_21# X VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
X0 VPWR VGND VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0.452 ps=4.52 w=0.87 l=2.89
X1 VGND VPWR VGND VNB sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0.286 ps=3.24 w=0.55 l=2.89
.ends

.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
X0 VPWR VGND VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0.452 ps=4.52 w=0.87 l=1.97
X1 VGND VPWR VGND VNB sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0.286 ps=3.24 w=0.55 l=1.97
.ends

.subckt sky130_fd_sc_hd__nor3b_1 A B C_N VGND VNB VPB VPWR Y
X0 VGND a_91_199# Y VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.221 ps=1.98 w=0.65 l=0.15
X1 Y B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X2 VPWR A a_245_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.146 pd=1.34 as=0.135 ps=1.27 w=1 l=0.15
X3 a_91_199# C_N VGND VNB sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.1 ps=0.985 w=0.42 l=0.15
X4 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.985 as=0.0878 ps=0.92 w=0.65 l=0.15
X5 a_245_297# B a_161_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6 a_91_199# C_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.146 ps=1.34 w=0.42 l=0.15
X7 a_161_297# a_91_199# Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.32 ps=2.64 w=1 l=0.15
.ends

.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
X0 VPWR VGND VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0.452 ps=4.52 w=0.87 l=1.05
X1 VGND VPWR VGND VNB sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0.286 ps=3.24 w=0.55 l=1.05
.ends

.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
X0 VPWR A a_110_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X5 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X6 a_110_47# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X7 a_110_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X8 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X9 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X10 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X11 a_110_47# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X12 VGND A a_110_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X13 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.0578 pd=0.695 as=0.0588 ps=0.7 w=0.42 l=0.15
X14 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X15 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X16 VGND A a_110_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X17 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.111 pd=1.37 as=0.0588 ps=0.7 w=0.42 l=0.15
X18 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.138 pd=1.27 as=0.14 ps=1.28 w=1 l=0.15
X19 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X20 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.138 ps=1.27 w=1 l=0.15
X21 a_110_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.111 ps=1.37 w=0.42 l=0.15
X22 VPWR A a_110_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X23 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X24 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X25 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X26 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X27 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X28 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X29 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X30 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X31 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X32 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X33 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X34 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X35 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X36 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X37 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X38 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X39 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0578 ps=0.695 w=0.42 l=0.15
.ends

.subckt sky130_ef_sc_hd__decap_12 VGND VPWR VPB VNB
X0 VPWR VGND VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0.452 ps=4.52 w=0.87 l=4.73
X1 VGND VPWR VGND VNB sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0.286 ps=3.24 w=0.55 l=4.73
.ends

.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
X0 VPWR A a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.162 pd=1.33 as=0.265 ps=2.53 w=1 l=0.15
X1 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2 VGND A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0683 pd=0.745 as=0.111 ps=1.37 w=0.42 l=0.15
X3 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.162 ps=1.33 w=1 l=0.15
X4 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0683 ps=0.745 w=0.42 l=0.15
X5 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
X0 VPWR a_75_212# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X1 a_75_212# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X2 a_75_212# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X3 VGND a_75_212# X VNB sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
.ends

.subckt sky130_fd_sc_hd__dlymetal6s2s_1 A VGND VNB VPB VPWR X
X0 a_558_47# a_381_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.141 ps=1.33 w=1 l=0.15
X1 VGND X a_381_47# VNB sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X2 a_841_47# a_664_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.141 ps=1.33 w=1 l=0.15
X3 VPWR A a_62_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.141 pd=1.33 as=0.109 ps=1.36 w=0.42 l=0.15
X4 VGND A a_62_47# VNB sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X5 a_558_47# a_381_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X6 X a_62_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.141 ps=1.33 w=1 l=0.15
X7 VPWR X a_381_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.141 pd=1.33 as=0.109 ps=1.36 w=0.42 l=0.15
X8 a_841_47# a_664_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X9 X a_62_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X10 VPWR a_558_47# a_664_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.141 pd=1.33 as=0.109 ps=1.36 w=0.42 l=0.15
X11 VGND a_558_47# a_664_47# VNB sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__dfrtp_1 CLK D RESET_B VGND VNB VPB VPWR Q
X0 a_1217_47# a_27_47# a_1108_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X1 a_805_47# a_761_289# a_639_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.14 ps=1.1 w=0.42 l=0.15
X2 a_1108_47# a_193_47# a_761_289# VNB sky130_fd_pr__nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X3 a_1283_21# a_1108_47# a_1462_47# VNB sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.064 ps=0.725 w=0.42 l=0.15
X4 a_651_413# a_27_47# a_543_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.116 pd=0.97 as=0.0724 ps=0.765 w=0.42 l=0.15
X5 VGND RESET_B a_805_47# VNB sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X6 Q a_1283_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.301 ps=2.66 w=1 l=0.15
X7 VPWR CLK a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X8 a_448_47# D VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.109 ps=1.36 w=0.42 l=0.15
X9 a_761_289# a_543_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.135 ps=1.15 w=0.64 l=0.15
X10 a_193_47# a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X11 a_1108_47# a_27_47# a_761_289# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.129 ps=1.18 w=0.42 l=0.15
X12 a_543_47# a_27_47# a_448_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X13 a_1462_47# RESET_B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.064 pd=0.725 as=0.125 ps=1.01 w=0.42 l=0.15
X14 a_543_47# a_193_47# a_448_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0724 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X15 a_448_47# D VGND VNB sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.221 ps=1.89 w=0.42 l=0.15
X16 VPWR a_1283_21# a_1270_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X17 VPWR a_1108_47# a_1283_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.113 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X18 a_1270_413# a_193_47# a_1108_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X19 a_193_47# a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X20 a_1283_21# RESET_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X21 VPWR a_761_289# a_651_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0703 pd=0.755 as=0.116 ps=0.97 w=0.42 l=0.15
X22 Q a_1283_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.209 ps=2.02 w=0.65 l=0.15
X23 a_639_47# a_193_47# a_543_47# VNB sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X24 VGND a_1283_21# a_1217_47# VNB sky130_fd_pr__nfet_01v8 ad=0.125 pd=1.01 as=0.0669 ps=0.75 w=0.42 l=0.15
X25 a_651_413# RESET_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0703 ps=0.755 w=0.42 l=0.15
X26 VGND CLK a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X27 a_761_289# a_543_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.129 pd=1.18 as=0.218 ps=2.2 w=0.84 l=0.15
.ends

.subckt sky130_fd_sc_hd__and2_1 A B VGND VNB VPB VPWR X
X0 VPWR B a_59_75# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.167 pd=1.39 as=0.0567 ps=0.69 w=0.42 l=0.15
X1 X a_59_75# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.475 pd=2.95 as=0.167 ps=1.39 w=1 l=0.15
X2 VGND B a_145_75# VNB sky130_fd_pr__nfet_01v8 ad=0.112 pd=1.04 as=0.0567 ps=0.69 w=0.42 l=0.15
X3 a_59_75# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.118 ps=1.4 w=0.42 l=0.15
X4 X a_59_75# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.112 ps=1.04 w=0.65 l=0.15
X5 a_145_75# A a_59_75# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.118 ps=1.4 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__dlygate4sd3_1 A VGND VNB VPB VPWR X
X0 VPWR A a_49_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X1 VGND a_285_47# a_391_47# VNB sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.5
X2 X a_391_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.141 ps=1.33 w=1 l=0.15
X3 VGND A a_49_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X4 VPWR a_285_47# a_391_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.141 pd=1.33 as=0.109 ps=1.36 w=0.42 l=0.5
X5 a_285_47# a_49_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.5
X6 a_285_47# a_49_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.5
X7 X a_391_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__nor2_2 A B VGND VNB VPB VPWR Y
X0 Y B a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1 Y B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X2 a_27_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X4 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.182 ps=1.86 w=0.65 l=0.15
X5 VGND B Y VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X6 VPWR A a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=2.56 w=1 l=0.15
X7 a_27_297# B Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
.ends

.subckt sky130_fd_sc_hd__o32a_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
X0 a_77_199# B2 a_227_47# VNB sky130_fd_pr__nfet_01v8 ad=0.133 pd=1.06 as=0.127 ps=1.04 w=0.65 l=0.15
X1 a_323_297# A2 a_227_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=1.39 as=0.165 ps=1.33 w=1 l=0.15
X2 a_227_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.135 ps=1.27 w=1 l=0.15
X3 a_227_47# B1 a_77_199# VNB sky130_fd_pr__nfet_01v8 ad=0.189 pd=1.88 as=0.133 ps=1.06 w=0.65 l=0.15
X4 VGND a_77_199# X VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5 VPWR B1 a_539_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.205 ps=1.41 w=1 l=0.15
X6 a_227_47# A3 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.127 pd=1.04 as=0.127 ps=1.04 w=0.65 l=0.15
X7 VPWR a_77_199# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.335 ps=2.67 w=1 l=0.15
X8 a_77_199# A3 a_323_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=1.39 as=0.195 ps=1.39 w=1 l=0.15
X9 VGND A2 a_227_47# VNB sky130_fd_pr__nfet_01v8 ad=0.127 pd=1.04 as=0.107 ps=0.98 w=0.65 l=0.15
X10 a_227_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.0878 ps=0.92 w=0.65 l=0.15
X11 a_539_297# B2 a_77_199# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=1.41 as=0.195 ps=1.39 w=1 l=0.15
.ends

.subckt scanchain data_out[0] data_out[1] data_out[2] data_out[3] data_out[4] data_out[5]
+ data_out[6] data_out[7] scan_out VDD GND
XPHY_EDGE_ROW_0_Left_12 GND GND VDD VDD sky130_fd_sc_hd__decap_3
X_66_ net1 _09_ _08_ GND GND VDD VDD _33_ sky130_fd_sc_hd__a21oi_1
X_49_ _11_ _18_ _19_ _20_ GND GND VDD VDD _02_ sky130_fd_sc_hd__o31a_1
Xoutput7 net7 GND GND VDD VDD data_out[1] sky130_fd_sc_hd__buf_2
X_65_ _11_ _30_ _31_ _32_ GND GND VDD VDD _06_ sky130_fd_sc_hd__o31a_1
XFILLER_0_9_39 GND GND VDD VDD sky130_fd_sc_hd__decap_3
X_48_ _12_ net1 net17 GND GND VDD VDD _20_ sky130_fd_sc_hd__or3_1
XPHY_EDGE_ROW_6_Right_6 GND GND VDD VDD sky130_fd_sc_hd__decap_3
Xoutput10 net10 GND GND VDD VDD data_out[4] sky130_fd_sc_hd__clkbuf_4
Xoutput8 net8 GND GND VDD VDD data_out[2] sky130_fd_sc_hd__buf_2
X_64_ net3 net1 net18 GND GND VDD VDD _32_ sky130_fd_sc_hd__or3_1
X_47_ _12_ _09_ net7 GND GND VDD VDD _19_ sky130_fd_sc_hd__o21a_1
XFILLER_0_9_3 GND GND VDD VDD sky130_fd_sc_hd__decap_8
Xoutput11 net11 GND GND VDD VDD data_out[5] sky130_fd_sc_hd__buf_2
Xoutput9 net9 GND GND VDD VDD data_out[3] sky130_fd_sc_hd__buf_2
X_63_ _12_ net5 net11 GND GND VDD VDD _31_ sky130_fd_sc_hd__o21a_1
XFILLER_0_10_22 GND GND VDD VDD sky130_fd_sc_hd__decap_6
X_46_ _08_ _09_ net9 GND GND VDD VDD _18_ sky130_fd_sc_hd__nor3b_1
XPHY_EDGE_ROW_4_Left_16 GND GND VDD VDD sky130_fd_sc_hd__decap_3
Xoutput12 net12 GND GND VDD VDD data_out[6] sky130_fd_sc_hd__buf_2
X_62_ _08_ _09_ net13 GND GND VDD VDD _30_ sky130_fd_sc_hd__nor3b_1
X_45_ _11_ _15_ _16_ _17_ GND GND VDD VDD _01_ sky130_fd_sc_hd__o31a_1
Xoutput13 net13 GND GND VDD VDD data_out[7] sky130_fd_sc_hd__clkbuf_4
X_61_ _11_ _27_ _28_ _29_ GND GND VDD VDD _05_ sky130_fd_sc_hd__o31a_1
X_44_ _12_ net1 net7 GND GND VDD VDD _17_ sky130_fd_sc_hd__or3_1
Xoutput14 net14 GND GND VDD VDD scan_out sky130_fd_sc_hd__clkbuf_4
X_60_ net3 net1 net11 GND GND VDD VDD _29_ sky130_fd_sc_hd__or3_1
X_43_ _08_ _09_ net6 GND GND VDD VDD _16_ sky130_fd_sc_hd__o21a_1
XPHY_EDGE_ROW_1_Right_1 GND GND VDD VDD sky130_fd_sc_hd__decap_3
X_42_ _08_ _09_ net8 GND GND VDD VDD _15_ sky130_fd_sc_hd__nor3b_1
XPHY_EDGE_ROW_11_Left_23 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_0_1_13 GND GND VDD VDD sky130_fd_sc_hd__decap_4
Xclkbuf_0_clk clkbuf_0_clk/A GND GND VDD VDD clknet_0_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_4_24 GND GND VDD VDD sky130_fd_sc_hd__decap_4
X_41_ _10_ _11_ _13_ _14_ GND GND VDD VDD _00_ sky130_fd_sc_hd__o31a_1
XFILLER_0_7_46 GND GND VDD VDD sky130_fd_sc_hd__decap_8
X_40_ _12_ net1 net6 GND GND VDD VDD _14_ sky130_fd_sc_hd__or3_1
XPHY_EDGE_ROW_5_Right_5 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_0_7_7 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_10_29 GND GND VDD VDD sky130_fd_sc_hd__decap_8
XFILLER_0_1_38 GND GND VDD VDD sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_11_Right_11 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_0_7_37 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_3_Left_15 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_0_5_6 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_0_11_41 GND VDD VDD GND sky130_ef_sc_hd__decap_12
Xinput1 input1/A GND GND VDD VDD net1 sky130_fd_sc_hd__buf_2
XPHY_EDGE_ROW_9_Right_9 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_0_11_53 GND GND VDD VDD sky130_fd_sc_hd__decap_3
Xinput2 reset GND GND VDD VDD net2 sky130_fd_sc_hd__clkbuf_4
Xinput3 input3/A GND GND VDD VDD net3 sky130_fd_sc_hd__clkbuf_2
XPHY_EDGE_ROW_7_Left_19 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_0_Right_0 GND GND VDD VDD sky130_fd_sc_hd__decap_3
Xinput4 input4/A GND GND VDD VDD net4 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_5_52 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_10_Left_22 GND GND VDD VDD sky130_fd_sc_hd__decap_3
X_76_ net13 GND GND VDD VDD net14 sky130_fd_sc_hd__clkbuf_1
Xinput5 input5/A GND GND VDD VDD net5 sky130_fd_sc_hd__dlymetal6s2s_1
X_59_ _12_ net5 net10 GND GND VDD VDD _28_ sky130_fd_sc_hd__o21a_1
X_58_ _08_ _09_ net12 GND GND VDD VDD _27_ sky130_fd_sc_hd__nor3b_1
X_75_ clknet_1_1__leaf_clk net16 net2 GND GND VDD VDD net13 sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_4_Right_4 GND GND VDD VDD sky130_fd_sc_hd__decap_3
X_74_ clknet_1_1__leaf_clk _06_ net2 GND GND VDD VDD net12 sky130_fd_sc_hd__dfrtp_1
X_57_ _11_ _24_ _25_ _26_ GND GND VDD VDD _04_ sky130_fd_sc_hd__o31a_1
X_73_ clknet_1_1__leaf_clk _05_ net2 GND GND VDD VDD net11 sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_2_Left_14 GND GND VDD VDD sky130_fd_sc_hd__decap_3
X_56_ net3 net1 net10 GND GND VDD VDD _26_ sky130_fd_sc_hd__or3_1
Xclkbuf_1_0__f_clk clknet_0_clk GND GND VDD VDD clknet_1_0__leaf_clk sky130_fd_sc_hd__clkbuf_16
X_39_ _12_ net4 GND GND VDD VDD _13_ sky130_fd_sc_hd__and2_1
X_72_ clknet_1_1__leaf_clk _04_ net2 GND GND VDD VDD net10 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_5_57 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_10_Right_10 GND GND VDD VDD sky130_fd_sc_hd__decap_3
X_55_ _12_ net5 net9 GND GND VDD VDD _25_ sky130_fd_sc_hd__o21a_1
X_38_ net3 GND GND VDD VDD _12_ sky130_fd_sc_hd__buf_2
Xhold1 net12 GND GND VDD VDD net15 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_8_Right_8 GND GND VDD VDD sky130_fd_sc_hd__decap_3
X_71_ clknet_1_0__leaf_clk _03_ net2 GND GND VDD VDD net9 sky130_fd_sc_hd__dfrtp_1
X_54_ _08_ _09_ net11 GND GND VDD VDD _24_ sky130_fd_sc_hd__nor3b_1
X_37_ net3 net1 GND GND VDD VDD _11_ sky130_fd_sc_hd__nor2_2
Xhold2 _07_ GND GND VDD VDD net16 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_8_25 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_0_11_29 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_70_ clknet_1_0__leaf_clk _02_ net2 GND GND VDD VDD net8 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_5_37 GND GND VDD VDD sky130_fd_sc_hd__decap_8
X_53_ _11_ _21_ _22_ _23_ GND GND VDD VDD _03_ sky130_fd_sc_hd__o31a_1
XPHY_EDGE_ROW_6_Left_18 GND GND VDD VDD sky130_fd_sc_hd__decap_3
X_36_ _08_ _09_ net7 GND GND VDD VDD _10_ sky130_fd_sc_hd__nor3b_1
XPHY_EDGE_ROW_9_Left_21 GND GND VDD VDD sky130_fd_sc_hd__decap_3
Xhold3 net8 GND GND VDD VDD net17 sky130_fd_sc_hd__dlygate4sd3_1
X_52_ _12_ net1 net9 GND GND VDD VDD _23_ sky130_fd_sc_hd__or3_1
X_35_ net5 GND GND VDD VDD _09_ sky130_fd_sc_hd__buf_2
Xhold4 net12 GND GND VDD VDD net18 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_10_9 GND GND VDD VDD sky130_fd_sc_hd__decap_8
X_51_ _12_ net5 net8 GND GND VDD VDD _22_ sky130_fd_sc_hd__o21a_1
XFILLER_0_2_29 GND GND VDD VDD sky130_fd_sc_hd__decap_4
X_34_ net3 GND GND VDD VDD _08_ sky130_fd_sc_hd__buf_2
XFILLER_0_5_18 GND GND VDD VDD sky130_fd_sc_hd__decap_8
XFILLER_0_6_61 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_0_6_3 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_50_ _08_ _09_ net10 GND GND VDD VDD _21_ sky130_fd_sc_hd__nor3b_1
Xclkbuf_1_1__f_clk clknet_0_clk GND GND VDD VDD clknet_1_1__leaf_clk sky130_fd_sc_hd__clkbuf_16
XPHY_EDGE_ROW_3_Right_3 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_0_3_52 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_1_Left_13 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_0_4_3 GND GND VDD VDD sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_7_Right_7 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_0_0_34 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_5_Left_17 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_0_0_46 GND GND VDD VDD sky130_fd_sc_hd__decap_8
XFILLER_0_0_57 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_8_Left_20 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_0_2_3 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_0_0_15 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_69_ clknet_1_0__leaf_clk _01_ net2 GND GND VDD VDD net7 sky130_fd_sc_hd__dfrtp_1
X_68_ clknet_1_0__leaf_clk _00_ net2 GND GND VDD VDD net6 sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_2_Right_2 GND GND VDD VDD sky130_fd_sc_hd__decap_3
X_67_ _08_ net1 net13 _33_ net15 GND GND VDD VDD _07_ sky130_fd_sc_hd__o32a_1
XFILLER_0_0_3 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_0_6_49 GND VDD VDD GND sky130_ef_sc_hd__decap_12
Xoutput6 net6 GND GND VDD VDD data_out[0] sky130_fd_sc_hd__clkbuf_4
C0 _09_ _08_ 2.33f
C1 _08_ VDD 2.09f
C2 VDD net1 5.95f
C3 VDD clknet_1_0__leaf_clk 2.53f
C4 VDD net9 2.27f
C5 VDD _12_ 2.83f
C6 VDD net2 2.2f
C7 VDD net6 2.06f
C8 net1 _12_ 2.74f
C9 VDD clknet_1_1__leaf_clk 2.8f
C10 _09_ VDD 2.97f
C11 net2 GND 5.94f
C12 net10 GND 3.07f
C13 net8 GND 2.48f
C14 _12_ GND 3.92f
C15 net1 GND 3.49f
C16 VDD GND 0.13p
C17 clknet_0_clk GND 2.69f
C18 _11_ GND 3.4f
C19 clkbuf_0_clk/A GND 3.74f
C20 _08_ GND 2.76f
C21 net3 GND 3.25f
C22 net7 GND 3.41f
.ends

.subckt sky130_fd_pr__nfet_01v8_HRDN5X a_n129_n130# a_n369_n42# a_543_64# a_63_n130#
+ a_159_64# a_n417_64# a_687_n42# a_303_n42# a_n561_n42# a_n321_n130# a_n749_n42#
+ a_639_n130# a_n81_n42# a_399_n42# a_n273_n42# a_15_n42# a_447_n130# a_n609_64# a_591_n42#
+ a_207_n42# a_n465_n42# a_351_64# a_255_n130# a_n33_64# a_n225_64# a_n705_n130# a_n177_n42#
+ a_n657_n42# a_495_n42# a_111_n42# a_n513_n130# VSUBS
X0 a_303_n42# a_255_n130# a_207_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X1 a_591_n42# a_543_64# a_495_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X2 a_207_n42# a_159_64# a_111_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X3 a_399_n42# a_351_64# a_303_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X4 a_495_n42# a_447_n130# a_399_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X5 a_687_n42# a_639_n130# a_591_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X6 a_n561_n42# a_n609_64# a_n657_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X7 a_n657_n42# a_n705_n130# a_n749_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X8 a_n465_n42# a_n513_n130# a_n561_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X9 a_n369_n42# a_n417_64# a_n465_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X10 a_15_n42# a_n33_64# a_n81_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X11 a_111_n42# a_63_n130# a_15_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X12 a_n273_n42# a_n321_n130# a_n369_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X13 a_n81_n42# a_n129_n130# a_n177_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X14 a_n177_n42# a_n225_64# a_n273_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
.ends

.subckt sky130_fd_pr__cap_mim_m3_1_MH6KF8 c1_n1046_n900# m3_n1086_n940# VSUBS
X0 c1_n1046_n900# m3_n1086_n940# sky130_fd_pr__cap_mim_m3_1 l=9 w=9
C0 m3_n1086_n940# c1_n1046_n900# 7.78f
C1 m3_n1086_n940# VSUBS 3.31f
.ends

.subckt nmos_dnw3 vin out1 out2 clk clkb vs VSUBS
X0 clkb clk vin vs sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.126 ps=1.44 w=0.42 l=0.15
X1 vin clkb clk vs sky130_fd_pr__nfet_01v8 ad=0.126 pd=1.44 as=0.13 ps=1.46 w=0.42 l=0.15
X2 out2 clk vin vs sky130_fd_pr__nfet_01v8 ad=1.65 pd=7.1 as=0.945 ps=3.63 w=3 l=1
X3 vin clkb out1 vs sky130_fd_pr__nfet_01v8 ad=0.945 pd=3.63 as=1.65 ps=7.1 w=3 l=1
C0 vs VSUBS 6.64f
.ends

.subckt sky130_fd_pr__pfet_01v8_FBZ64Q a_n81_n126# a_399_n126# a_351_n223# a_n417_n223#
+ a_207_n126# a_n225_n223# a_n461_n126# a_n369_n126# a_63_157# a_303_n126# a_255_157#
+ a_n33_n223# a_15_n126# a_n177_n126# a_n129_157# a_111_n126# w_n497_n226# a_n273_n126#
+ a_159_n223# a_n321_157# VSUBS
X0 a_n273_n126# a_n321_157# a_n369_n126# w_n497_n226# sky130_fd_pr__pfet_01v8 ad=0.208 pd=1.59 as=0.208 ps=1.59 w=1.26 l=0.15
X1 a_207_n126# a_159_n223# a_111_n126# w_n497_n226# sky130_fd_pr__pfet_01v8 ad=0.208 pd=1.59 as=0.208 ps=1.59 w=1.26 l=0.15
X2 a_n177_n126# a_n225_n223# a_n273_n126# w_n497_n226# sky130_fd_pr__pfet_01v8 ad=0.208 pd=1.59 as=0.208 ps=1.59 w=1.26 l=0.15
X3 a_111_n126# a_63_157# a_15_n126# w_n497_n226# sky130_fd_pr__pfet_01v8 ad=0.208 pd=1.59 as=0.208 ps=1.59 w=1.26 l=0.15
X4 a_399_n126# a_351_n223# a_303_n126# w_n497_n226# sky130_fd_pr__pfet_01v8 ad=0.391 pd=3.14 as=0.208 ps=1.59 w=1.26 l=0.15
X5 a_n81_n126# a_n129_157# a_n177_n126# w_n497_n226# sky130_fd_pr__pfet_01v8 ad=0.208 pd=1.59 as=0.208 ps=1.59 w=1.26 l=0.15
X6 a_15_n126# a_n33_n223# a_n81_n126# w_n497_n226# sky130_fd_pr__pfet_01v8 ad=0.208 pd=1.59 as=0.208 ps=1.59 w=1.26 l=0.15
X7 a_n369_n126# a_n417_n223# a_n461_n126# w_n497_n226# sky130_fd_pr__pfet_01v8 ad=0.208 pd=1.59 as=0.391 ps=3.14 w=1.26 l=0.15
X8 a_303_n126# a_255_157# a_207_n126# w_n497_n226# sky130_fd_pr__pfet_01v8 ad=0.208 pd=1.59 as=0.208 ps=1.59 w=1.26 l=0.15
.ends

.subckt sky130_fd_pr__nfet_01v8_5ACVEW a_n129_n130# a_63_n130# a_n81_n42# a_15_n42#
+ a_n173_n42# a_n33_64# a_111_n42# VSUBS
X0 a_15_n42# a_n33_64# a_n81_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X1 a_111_n42# a_63_n130# a_15_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X2 a_n81_n42# a_n129_n130# a_n173_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
.ends

.subckt sky130_fd_pr__nfet_01v8_NJGLN5 a_n129_n130# a_n369_n42# a_1215_n130# a_543_64#
+ a_63_n130# a_159_64# a_n1089_n130# a_n849_n42# a_n417_64# a_n801_64# a_687_n42#
+ a_303_n42# a_1167_n42# a_n561_n42# a_n321_n130# a_n1041_n42# a_639_n130# a_n1185_64#
+ a_1023_n130# a_n1281_n130# a_n81_n42# a_399_n42# a_879_n42# a_n273_n42# a_735_64#
+ a_n753_n42# a_15_n42# a_n897_n130# a_n1233_n42# a_831_n130# a_447_n130# a_n609_64#
+ a_1071_n42# a_591_n42# a_1119_64# a_n993_64# a_207_n42# a_n465_n42# a_n945_n42#
+ a_351_64# a_783_n42# a_255_n130# a_n33_64# a_n225_64# a_n705_n130# a_1263_n42# a_927_64#
+ a_n177_n42# a_n657_n42# a_n1325_n42# a_n1137_n42# a_495_n42# a_111_n42# a_975_n42#
+ a_n513_n130# VSUBS
X0 a_303_n42# a_255_n130# a_207_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X1 a_591_n42# a_543_64# a_495_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X2 a_207_n42# a_159_64# a_111_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X3 a_399_n42# a_351_64# a_303_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X4 a_495_n42# a_447_n130# a_399_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X5 a_687_n42# a_639_n130# a_591_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X6 a_783_n42# a_735_64# a_687_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X7 a_975_n42# a_927_64# a_879_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X8 a_n1041_n42# a_n1089_n130# a_n1137_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X9 a_879_n42# a_831_n130# a_783_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X10 a_n1233_n42# a_n1281_n130# a_n1325_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X11 a_n1137_n42# a_n1185_64# a_n1233_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X12 a_n561_n42# a_n609_64# a_n657_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X13 a_1071_n42# a_1023_n130# a_975_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X14 a_1263_n42# a_1215_n130# a_1167_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X15 a_n945_n42# a_n993_64# a_n1041_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X16 a_n753_n42# a_n801_64# a_n849_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X17 a_n657_n42# a_n705_n130# a_n753_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X18 a_n465_n42# a_n513_n130# a_n561_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X19 a_n369_n42# a_n417_64# a_n465_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X20 a_1167_n42# a_1119_64# a_1071_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X21 a_n849_n42# a_n897_n130# a_n945_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X22 a_15_n42# a_n33_64# a_n81_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X23 a_111_n42# a_63_n130# a_15_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X24 a_n273_n42# a_n321_n130# a_n369_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X25 a_n81_n42# a_n129_n130# a_n177_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X26 a_n177_n42# a_n225_64# a_n273_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
.ends

.subckt sky130_fd_pr__pfet_01v8_VR4B8J a_1119_157# a_783_n126# a_n81_n126# a_n849_n126#
+ a_399_n126# a_n1041_n126# a_351_157# a_495_n126# a_n945_n126# a_n33_157# a_n129_n223#
+ a_n513_n223# a_1215_n223# a_63_n223# a_n1089_n223# a_n225_157# a_591_n126# a_n657_n126#
+ a_207_n126# a_543_157# a_n1325_n126# a_n369_n126# a_n753_n126# a_n321_n223# a_303_n126#
+ a_1023_n223# a_639_n223# a_n1281_n223# a_n417_157# a_n465_n126# a_1167_n126# a_735_157#
+ a_15_n126# a_n561_n126# a_n993_157# a_n177_n126# a_n897_n223# w_n1361_n226# a_1263_n126#
+ a_879_n126# a_111_n126# a_831_n223# a_n609_157# a_447_n223# a_n273_n126# a_n1137_n126#
+ a_975_n126# a_927_157# a_n1185_157# a_n1233_n126# a_n801_157# a_1071_n126# a_687_n126#
+ a_255_n223# a_n705_n223# a_159_157# VSUBS
X0 a_n273_n126# a_n321_n223# a_n369_n126# w_n1361_n226# sky130_fd_pr__pfet_01v8 ad=0.208 pd=1.59 as=0.208 ps=1.59 w=1.26 l=0.15
X1 a_n1233_n126# a_n1281_n223# a_n1325_n126# w_n1361_n226# sky130_fd_pr__pfet_01v8 ad=0.208 pd=1.59 as=0.391 ps=3.14 w=1.26 l=0.15
X2 a_591_n126# a_543_157# a_495_n126# w_n1361_n226# sky130_fd_pr__pfet_01v8 ad=0.208 pd=1.59 as=0.208 ps=1.59 w=1.26 l=0.15
X3 a_n849_n126# a_n897_n223# a_n945_n126# w_n1361_n226# sky130_fd_pr__pfet_01v8 ad=0.208 pd=1.59 as=0.208 ps=1.59 w=1.26 l=0.15
X4 a_207_n126# a_159_157# a_111_n126# w_n1361_n226# sky130_fd_pr__pfet_01v8 ad=0.208 pd=1.59 as=0.208 ps=1.59 w=1.26 l=0.15
X5 a_n177_n126# a_n225_157# a_n273_n126# w_n1361_n226# sky130_fd_pr__pfet_01v8 ad=0.208 pd=1.59 as=0.208 ps=1.59 w=1.26 l=0.15
X6 a_n1137_n126# a_n1185_157# a_n1233_n126# w_n1361_n226# sky130_fd_pr__pfet_01v8 ad=0.208 pd=1.59 as=0.208 ps=1.59 w=1.26 l=0.15
X7 a_495_n126# a_447_n223# a_399_n126# w_n1361_n226# sky130_fd_pr__pfet_01v8 ad=0.208 pd=1.59 as=0.208 ps=1.59 w=1.26 l=0.15
X8 a_n561_n126# a_n609_157# a_n657_n126# w_n1361_n226# sky130_fd_pr__pfet_01v8 ad=0.208 pd=1.59 as=0.208 ps=1.59 w=1.26 l=0.15
X9 a_111_n126# a_63_n223# a_15_n126# w_n1361_n226# sky130_fd_pr__pfet_01v8 ad=0.208 pd=1.59 as=0.208 ps=1.59 w=1.26 l=0.15
X10 a_783_n126# a_735_157# a_687_n126# w_n1361_n226# sky130_fd_pr__pfet_01v8 ad=0.208 pd=1.59 as=0.208 ps=1.59 w=1.26 l=0.15
X11 a_1071_n126# a_1023_n223# a_975_n126# w_n1361_n226# sky130_fd_pr__pfet_01v8 ad=0.208 pd=1.59 as=0.208 ps=1.59 w=1.26 l=0.15
X12 a_399_n126# a_351_157# a_303_n126# w_n1361_n226# sky130_fd_pr__pfet_01v8 ad=0.208 pd=1.59 as=0.208 ps=1.59 w=1.26 l=0.15
X13 a_n465_n126# a_n513_n223# a_n561_n126# w_n1361_n226# sky130_fd_pr__pfet_01v8 ad=0.208 pd=1.59 as=0.208 ps=1.59 w=1.26 l=0.15
X14 a_687_n126# a_639_n223# a_591_n126# w_n1361_n226# sky130_fd_pr__pfet_01v8 ad=0.208 pd=1.59 as=0.208 ps=1.59 w=1.26 l=0.15
X15 a_n753_n126# a_n801_157# a_n849_n126# w_n1361_n226# sky130_fd_pr__pfet_01v8 ad=0.208 pd=1.59 as=0.208 ps=1.59 w=1.26 l=0.15
X16 a_975_n126# a_927_157# a_879_n126# w_n1361_n226# sky130_fd_pr__pfet_01v8 ad=0.208 pd=1.59 as=0.208 ps=1.59 w=1.26 l=0.15
X17 a_n81_n126# a_n129_n223# a_n177_n126# w_n1361_n226# sky130_fd_pr__pfet_01v8 ad=0.208 pd=1.59 as=0.208 ps=1.59 w=1.26 l=0.15
X18 a_15_n126# a_n33_157# a_n81_n126# w_n1361_n226# sky130_fd_pr__pfet_01v8 ad=0.208 pd=1.59 as=0.208 ps=1.59 w=1.26 l=0.15
X19 a_1263_n126# a_1215_n223# a_1167_n126# w_n1361_n226# sky130_fd_pr__pfet_01v8 ad=0.391 pd=3.14 as=0.208 ps=1.59 w=1.26 l=0.15
X20 a_n1041_n126# a_n1089_n223# a_n1137_n126# w_n1361_n226# sky130_fd_pr__pfet_01v8 ad=0.208 pd=1.59 as=0.208 ps=1.59 w=1.26 l=0.15
X21 a_n369_n126# a_n417_157# a_n465_n126# w_n1361_n226# sky130_fd_pr__pfet_01v8 ad=0.208 pd=1.59 as=0.208 ps=1.59 w=1.26 l=0.15
X22 a_n657_n126# a_n705_n223# a_n753_n126# w_n1361_n226# sky130_fd_pr__pfet_01v8 ad=0.208 pd=1.59 as=0.208 ps=1.59 w=1.26 l=0.15
X23 a_879_n126# a_831_n223# a_783_n126# w_n1361_n226# sky130_fd_pr__pfet_01v8 ad=0.208 pd=1.59 as=0.208 ps=1.59 w=1.26 l=0.15
X24 a_n945_n126# a_n993_157# a_n1041_n126# w_n1361_n226# sky130_fd_pr__pfet_01v8 ad=0.208 pd=1.59 as=0.208 ps=1.59 w=1.26 l=0.15
X25 a_1167_n126# a_1119_157# a_1071_n126# w_n1361_n226# sky130_fd_pr__pfet_01v8 ad=0.208 pd=1.59 as=0.208 ps=1.59 w=1.26 l=0.15
X26 a_303_n126# a_255_n223# a_207_n126# w_n1361_n226# sky130_fd_pr__pfet_01v8 ad=0.208 pd=1.59 as=0.208 ps=1.59 w=1.26 l=0.15
C0 w_n1361_n226# VSUBS 3.67f
.ends

.subckt inverter_27x m1_n804_1398# m1_540_1398# m1_156_1398# m1_n36_1398# m1_732_1398#
+ m1_n1102_1398# m1_348_1398# m1_n1188_1398# m1_n996_1398# m1_n228_1398# m1_n1188_1912#
+ m1_924_1398# m1_1309_1398# a_n1158_1658# m1_n420_1398# m1_1116_1398# w_1358_2036#
+ m1_n612_1398# VSUBS
Xsky130_fd_pr__nfet_01v8_NJGLN5_1 a_n1158_1658# m1_n228_1398# a_n1158_1658# a_n1158_1658#
+ a_n1158_1658# a_n1158_1658# a_n1158_1658# m1_n1102_1398# a_n1158_1658# a_n1158_1658#
+ m1_n1102_1398# m1_n1102_1398# m1_1309_1398# m1_n420_1398# a_n1158_1658# m1_n1102_1398#
+ a_n1158_1658# a_n1158_1658# a_n1158_1658# a_n1158_1658# m1_n1102_1398# m1_540_1398#
+ m1_n1102_1398# m1_n1102_1398# a_n1158_1658# m1_n612_1398# m1_156_1398# a_n1158_1658#
+ m1_n1102_1398# a_n1158_1658# a_n1158_1658# a_n1158_1658# m1_n1102_1398# m1_732_1398#
+ a_n1158_1658# a_n1158_1658# m1_348_1398# m1_n1102_1398# m1_n804_1398# a_n1158_1658#
+ m1_924_1398# a_n1158_1658# a_n1158_1658# a_n1158_1658# a_n1158_1658# m1_n1102_1398#
+ a_n1158_1658# m1_n36_1398# m1_n1102_1398# m1_n1188_1398# m1_n996_1398# m1_n1102_1398#
+ m1_n1102_1398# m1_1116_1398# a_n1158_1658# VSUBS sky130_fd_pr__nfet_01v8_NJGLN5
Xsky130_fd_pr__pfet_01v8_VR4B8J_1 a_n1158_1658# m1_n1188_1912# m1_1309_1398# m1_1309_1398#
+ m1_n1188_1912# m1_1309_1398# a_n1158_1658# m1_1309_1398# m1_n1188_1912# a_n1158_1658#
+ a_n1158_1658# a_n1158_1658# a_n1158_1658# a_n1158_1658# a_n1158_1658# a_n1158_1658#
+ m1_n1188_1912# m1_1309_1398# m1_n1188_1912# a_n1158_1658# m1_n1188_1912# m1_n1188_1912#
+ m1_n1188_1912# a_n1158_1658# m1_1309_1398# a_n1158_1658# a_n1158_1658# a_n1158_1658#
+ a_n1158_1658# m1_1309_1398# m1_n1188_1912# a_n1158_1658# m1_n1188_1912# m1_n1188_1912#
+ a_n1158_1658# m1_n1188_1912# a_n1158_1658# w_1358_2036# m1_1309_1398# m1_1309_1398#
+ m1_1309_1398# a_n1158_1658# a_n1158_1658# a_n1158_1658# m1_1309_1398# m1_n1188_1912#
+ m1_n1188_1912# a_n1158_1658# a_n1158_1658# m1_1309_1398# a_n1158_1658# m1_1309_1398#
+ m1_1309_1398# a_n1158_1658# a_n1158_1658# a_n1158_1658# VSUBS sky130_fd_pr__pfet_01v8_VR4B8J
C0 a_n1158_1658# VSUBS 6.39f
C1 w_1358_2036# VSUBS 3.69f
.ends

.subckt sky130_fd_pr__nfet_01v8_KMMFCM a_15_n42# a_n15_n68# a_n73_n42# VSUBS
X0 a_15_n42# a_n15_n68# a_n73_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
.ends

.subckt sky130_fd_pr__pfet_01v8_29EZRJ a_n73_n126# w_n109_n188# a_15_n126# a_n15_n152#
+ VSUBS
X0 a_15_n126# a_n15_n152# a_n73_n126# w_n109_n188# sky130_fd_pr__pfet_01v8 ad=0.365 pd=3.1 as=0.365 ps=3.1 w=1.26 l=0.15
.ends

.subckt sky130_fd_pr__pfet_01v8_FL984Q a_n81_n126# a_n33_157# a_n129_n223# a_63_n223#
+ a_n173_n126# a_15_n126# a_111_n126# w_n209_n226# VSUBS
X0 a_111_n126# a_63_n223# a_15_n126# w_n209_n226# sky130_fd_pr__pfet_01v8 ad=0.391 pd=3.14 as=0.208 ps=1.59 w=1.26 l=0.15
X1 a_n81_n126# a_n129_n223# a_n173_n126# w_n209_n226# sky130_fd_pr__pfet_01v8 ad=0.208 pd=1.59 as=0.391 ps=3.14 w=1.26 l=0.15
X2 a_15_n126# a_n33_157# a_n81_n126# w_n209_n226# sky130_fd_pr__pfet_01v8 ad=0.208 pd=1.59 as=0.208 ps=1.59 w=1.26 l=0.15
.ends

.subckt sky130_fd_pr__pfet_01v8_FXZ64Q a_n73_n126# w_n109_n188# a_15_n126# a_n15_n152#
+ VSUBS
X0 a_15_n126# a_n15_n152# a_n73_n126# w_n109_n188# sky130_fd_pr__pfet_01v8 ad=0.365 pd=3.1 as=0.365 ps=3.1 w=1.26 l=0.15
.ends

.subckt sky130_fd_pr__nfet_01v8_D4CDWR a_n369_n42# a_n225_n130# a_303_n42# a_n81_n42#
+ a_399_n42# a_n33_n130# a_n273_n42# a_n461_n42# a_15_n42# a_n321_64# a_207_n42# a_159_n130#
+ a_n177_n42# a_351_n130# a_255_64# a_n417_n130# a_111_n42# a_n129_64# a_63_64# VSUBS
X0 a_303_n42# a_255_64# a_207_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X1 a_207_n42# a_159_n130# a_111_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X2 a_399_n42# a_351_n130# a_303_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X3 a_n369_n42# a_n417_n130# a_n461_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X4 a_15_n42# a_n33_n130# a_n81_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X5 a_111_n42# a_63_64# a_15_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X6 a_n273_n42# a_n321_64# a_n369_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X7 a_n81_n42# a_n129_64# a_n177_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X8 a_n177_n42# a_n225_n130# a_n273_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
.ends

.subckt sky130_fd_pr__nfet_01v8_DQBD8A a_15_n42# a_n15_n68# a_n73_n42# VSUBS
X0 a_15_n42# a_n15_n68# a_n73_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
.ends

.subckt clock clk_in vdd gnd clk clkb
Xsky130_fd_pr__pfet_01v8_FBZ64Q_0 vdd a_3246_118# a_2402_572# a_2402_572# a_3246_118#
+ a_2402_572# vdd a_3246_118# a_2402_572# vdd a_2402_572# a_2402_572# a_3246_118#
+ a_3246_118# a_2402_572# vdd vdd vdd a_2402_572# a_2402_572# gnd sky130_fd_pr__pfet_01v8_FBZ64Q
Xsky130_fd_pr__nfet_01v8_5ACVEW_0 a_344_n986# a_344_n986# a_2402_572# gnd gnd a_344_n986#
+ a_2402_572# gnd sky130_fd_pr__nfet_01v8_5ACVEW
Xinverter_27x_0 clk clk clk clk clk gnd clk clk clk clk vdd clk clk a_3246_118# clk
+ clk vdd clk gnd inverter_27x
Xsky130_fd_pr__nfet_01v8_KMMFCM_0 a_134_122# clk_in gnd gnd sky130_fd_pr__nfet_01v8_KMMFCM
Xsky130_fd_pr__nfet_01v8_KMMFCM_1 a_416_120# a_344_102# sky130_fd_pr__nfet_01v8_KMMFCM_2/a_15_n42#
+ gnd sky130_fd_pr__nfet_01v8_KMMFCM
Xsky130_fd_pr__nfet_01v8_KMMFCM_2 sky130_fd_pr__nfet_01v8_KMMFCM_2/a_15_n42# a_134_122#
+ gnd gnd sky130_fd_pr__nfet_01v8_KMMFCM
Xsky130_fd_pr__pfet_01v8_29EZRJ_0 vdd vdd a_134_122# clk_in gnd sky130_fd_pr__pfet_01v8_29EZRJ
Xsky130_fd_pr__pfet_01v8_FL984Q_0 a_2402_572# a_344_n986# a_344_n986# a_344_n986#
+ vdd vdd a_2402_572# vdd gnd sky130_fd_pr__pfet_01v8_FL984Q
Xsky130_fd_pr__pfet_01v8_FXZ64Q_0 vdd vdd a_1230_122# m1_998_498# gnd sky130_fd_pr__pfet_01v8_FXZ64Q
Xsky130_fd_pr__pfet_01v8_29EZRJ_1 a_416_120# vdd vdd a_344_102# gnd sky130_fd_pr__pfet_01v8_29EZRJ
Xsky130_fd_pr__pfet_01v8_FXZ64Q_1 vdd vdd a_1430_122# a_1230_122# gnd sky130_fd_pr__pfet_01v8_FXZ64Q
Xsky130_fd_pr__pfet_01v8_29EZRJ_2 vdd vdd a_416_120# a_134_122# gnd sky130_fd_pr__pfet_01v8_29EZRJ
Xsky130_fd_pr__pfet_01v8_FXZ64Q_2 vdd vdd a_344_n986# a_1430_122# gnd sky130_fd_pr__pfet_01v8_FXZ64Q
Xsky130_fd_pr__pfet_01v8_29EZRJ_3 vdd vdd m1_998_498# a_786_n2# gnd sky130_fd_pr__pfet_01v8_29EZRJ
Xsky130_fd_pr__nfet_01v8_D4CDWR_0 a_3246_118# a_2402_572# gnd gnd a_3246_118# a_2402_572#
+ gnd gnd a_3246_118# a_2402_572# a_3246_118# a_2402_572# a_3246_118# a_2402_572#
+ a_2402_572# a_2402_572# gnd a_2402_572# a_2402_572# gnd sky130_fd_pr__nfet_01v8_D4CDWR
Xsky130_fd_pr__nfet_01v8_DQBD8A_0 m1_998_498# a_786_n2# gnd gnd sky130_fd_pr__nfet_01v8_DQBD8A
Xsky130_fd_pr__nfet_01v8_DQBD8A_1 a_1230_122# m1_998_498# gnd gnd sky130_fd_pr__nfet_01v8_DQBD8A
Xsky130_fd_pr__nfet_01v8_DQBD8A_2 a_1430_122# a_1230_122# gnd gnd sky130_fd_pr__nfet_01v8_DQBD8A
Xsky130_fd_pr__nfet_01v8_DQBD8A_3 a_344_n986# a_1430_122# gnd gnd sky130_fd_pr__nfet_01v8_DQBD8A
X0 gnd a_2432_n962# clkb gnd sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X1 vdd a_2432_n962# clkb vdd sky130_fd_pr__pfet_01v8 ad=0.208 pd=1.59 as=0.208 ps=1.59 w=1.26 l=0.15
X2 vdd a_2020_n482# a_2432_n962# vdd sky130_fd_pr__pfet_01v8 ad=0.208 pd=1.59 as=0.208 ps=1.59 w=1.26 l=0.15
X3 clkb a_2432_n962# gnd gnd sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X4 vdd a_344_102# a_2020_n482# vdd sky130_fd_pr__pfet_01v8 ad=0.208 pd=1.59 as=0.208 ps=1.59 w=1.26 l=0.15
X5 gnd a_2432_n962# clkb gnd sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X6 vdd a_2432_n962# clkb vdd sky130_fd_pr__pfet_01v8 ad=0.208 pd=1.59 as=0.208 ps=1.59 w=1.26 l=0.15
X7 clkb a_2432_n962# gnd gnd sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X8 a_2020_n482# a_344_102# gnd gnd sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X9 a_786_n912# a_586_n912# vdd vdd sky130_fd_pr__pfet_01v8 ad=0.365 pd=3.1 as=0.365 ps=3.1 w=1.26 l=0.15
X10 vdd a_2432_n962# clkb vdd sky130_fd_pr__pfet_01v8 ad=0.208 pd=1.59 as=0.208 ps=1.59 w=1.26 l=0.15
X11 a_2432_n962# a_2020_n482# vdd vdd sky130_fd_pr__pfet_01v8 ad=0.208 pd=1.59 as=0.208 ps=1.59 w=1.26 l=0.15
X12 clkb a_2432_n962# vdd vdd sky130_fd_pr__pfet_01v8 ad=0.208 pd=1.59 as=0.208 ps=1.59 w=1.26 l=0.15
X13 clkb a_2432_n962# gnd gnd sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X14 gnd a_2020_n482# a_2432_n962# gnd sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X15 clkb a_2432_n962# gnd gnd sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X16 clkb a_2432_n962# vdd vdd sky130_fd_pr__pfet_01v8 ad=0.208 pd=1.59 as=0.208 ps=1.59 w=1.26 l=0.15
X17 gnd a_2432_n962# clkb gnd sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X18 gnd a_2020_n482# a_2432_n962# gnd sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X19 vdd a_2432_n962# clkb vdd sky130_fd_pr__pfet_01v8 ad=0.208 pd=1.59 as=0.208 ps=1.59 w=1.26 l=0.15
X20 a_286_n478# clk_in gnd gnd sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0.122 ps=1.42 w=0.42 l=0.15
X21 clkb a_2432_n962# vdd vdd sky130_fd_pr__pfet_01v8 ad=0.208 pd=1.59 as=0.208 ps=1.59 w=1.26 l=0.15
X22 gnd a_2432_n962# clkb gnd sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X23 a_2432_n962# a_2020_n482# vdd vdd sky130_fd_pr__pfet_01v8 ad=0.208 pd=1.59 as=0.391 ps=3.14 w=1.26 l=0.15
X24 clkb a_2432_n962# gnd gnd sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X25 a_2432_n962# a_2020_n482# gnd gnd sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X26 a_586_n2# a_416_120# gnd gnd sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X27 clkb a_2432_n962# vdd vdd sky130_fd_pr__pfet_01v8 ad=0.208 pd=1.59 as=0.208 ps=1.59 w=1.26 l=0.15
X28 gnd a_2432_n962# clkb gnd sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X29 a_2432_n962# a_2020_n482# vdd vdd sky130_fd_pr__pfet_01v8 ad=0.391 pd=3.14 as=0.208 ps=1.59 w=1.26 l=0.15
X30 a_786_n912# a_586_n912# gnd gnd sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X31 clkb a_2432_n962# vdd vdd sky130_fd_pr__pfet_01v8 ad=0.208 pd=1.59 as=0.208 ps=1.59 w=1.26 l=0.15
X32 gnd a_2432_n962# clkb gnd sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X33 vdd a_344_n986# a_286_n960# vdd sky130_fd_pr__pfet_01v8 ad=0.365 pd=3.1 as=0.183 ps=1.55 w=1.26 l=0.15
X34 a_344_102# a_1394_n918# vdd vdd sky130_fd_pr__pfet_01v8 ad=0.365 pd=3.1 as=0.365 ps=3.1 w=1.26 l=0.15
X35 a_992_n918# a_786_n912# vdd vdd sky130_fd_pr__pfet_01v8 ad=0.365 pd=3.1 as=0.365 ps=3.1 w=1.26 l=0.15
X36 a_1192_n918# a_992_n918# gnd gnd sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X37 vdd a_2432_n962# clkb vdd sky130_fd_pr__pfet_01v8 ad=0.208 pd=1.59 as=0.208 ps=1.59 w=1.26 l=0.15
X38 a_2432_n962# a_2020_n482# vdd vdd sky130_fd_pr__pfet_01v8 ad=0.208 pd=1.59 as=0.208 ps=1.59 w=1.26 l=0.15
X39 gnd a_2432_n962# clkb gnd sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X40 a_2432_n962# a_2020_n482# gnd gnd sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X41 a_1394_n918# a_1192_n918# gnd gnd sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X42 vdd a_2432_n962# clkb vdd sky130_fd_pr__pfet_01v8 ad=0.208 pd=1.59 as=0.208 ps=1.59 w=1.26 l=0.15
X43 clkb a_2432_n962# gnd gnd sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X44 clkb a_2432_n962# gnd gnd sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X45 clkb a_2432_n962# vdd vdd sky130_fd_pr__pfet_01v8 ad=0.208 pd=1.59 as=0.208 ps=1.59 w=1.26 l=0.15
X46 gnd a_2020_n482# a_2432_n962# gnd sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X47 vdd a_2432_n962# clkb vdd sky130_fd_pr__pfet_01v8 ad=0.208 pd=1.59 as=0.208 ps=1.59 w=1.26 l=0.15
X48 vdd a_2020_n482# a_2432_n962# vdd sky130_fd_pr__pfet_01v8 ad=0.208 pd=1.59 as=0.208 ps=1.59 w=1.26 l=0.15
X49 gnd a_2432_n962# clkb gnd sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X50 a_2020_n482# a_344_102# vdd vdd sky130_fd_pr__pfet_01v8 ad=0.391 pd=3.14 as=0.208 ps=1.59 w=1.26 l=0.15
X51 vdd a_2432_n962# clkb vdd sky130_fd_pr__pfet_01v8 ad=0.208 pd=1.59 as=0.208 ps=1.59 w=1.26 l=0.15
X52 clkb a_2432_n962# gnd gnd sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X53 a_586_n912# a_286_n960# vdd vdd sky130_fd_pr__pfet_01v8 ad=0.365 pd=3.1 as=0.365 ps=3.1 w=1.26 l=0.15
X54 vdd a_2020_n482# a_2432_n962# vdd sky130_fd_pr__pfet_01v8 ad=0.208 pd=1.59 as=0.208 ps=1.59 w=1.26 l=0.15
X55 a_586_n2# a_416_120# vdd vdd sky130_fd_pr__pfet_01v8 ad=0.365 pd=3.1 as=0.365 ps=3.1 w=1.26 l=0.15
X56 clkb a_2432_n962# vdd vdd sky130_fd_pr__pfet_01v8 ad=0.208 pd=1.59 as=0.391 ps=3.14 w=1.26 l=0.15
X57 clkb a_2432_n962# vdd vdd sky130_fd_pr__pfet_01v8 ad=0.208 pd=1.59 as=0.208 ps=1.59 w=1.26 l=0.15
X58 vdd a_2432_n962# clkb vdd sky130_fd_pr__pfet_01v8 ad=0.208 pd=1.59 as=0.208 ps=1.59 w=1.26 l=0.15
X59 clkb a_2432_n962# gnd gnd sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X60 gnd a_2432_n962# clkb gnd sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X61 gnd a_2020_n482# a_2432_n962# gnd sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X62 clkb a_2432_n962# vdd vdd sky130_fd_pr__pfet_01v8 ad=0.208 pd=1.59 as=0.208 ps=1.59 w=1.26 l=0.15
X63 gnd a_2432_n962# clkb gnd sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X64 clkb a_2432_n962# gnd gnd sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X65 clkb a_2432_n962# vdd vdd sky130_fd_pr__pfet_01v8 ad=0.208 pd=1.59 as=0.208 ps=1.59 w=1.26 l=0.15
X66 a_2020_n482# a_344_102# gnd gnd sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X67 vdd a_2432_n962# clkb vdd sky130_fd_pr__pfet_01v8 ad=0.208 pd=1.59 as=0.208 ps=1.59 w=1.26 l=0.15
X68 gnd a_2432_n962# clkb gnd sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X69 a_2432_n962# a_2020_n482# gnd gnd sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X70 gnd a_2432_n962# clkb gnd sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X71 a_786_n2# a_586_n2# gnd gnd sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X72 clkb a_2432_n962# gnd gnd sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X73 a_286_n960# clk_in vdd vdd sky130_fd_pr__pfet_01v8 ad=0.183 pd=1.55 as=0.365 ps=3.1 w=1.26 l=0.15
X74 clkb a_2432_n962# vdd vdd sky130_fd_pr__pfet_01v8 ad=0.208 pd=1.59 as=0.208 ps=1.59 w=1.26 l=0.15
X75 a_286_n960# a_344_n986# a_286_n478# gnd sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0609 ps=0.71 w=0.42 l=0.15
X76 a_2432_n962# a_2020_n482# vdd vdd sky130_fd_pr__pfet_01v8 ad=0.208 pd=1.59 as=0.208 ps=1.59 w=1.26 l=0.15
X77 a_586_n912# a_286_n960# gnd gnd sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X78 a_1394_n918# a_1192_n918# vdd vdd sky130_fd_pr__pfet_01v8 ad=0.365 pd=3.1 as=0.365 ps=3.1 w=1.26 l=0.15
X79 a_1192_n918# a_992_n918# vdd vdd sky130_fd_pr__pfet_01v8 ad=0.365 pd=3.1 as=0.365 ps=3.1 w=1.26 l=0.15
X80 gnd a_2432_n962# clkb gnd sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X81 a_2432_n962# a_2020_n482# gnd gnd sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X82 vdd a_2432_n962# clkb vdd sky130_fd_pr__pfet_01v8 ad=0.208 pd=1.59 as=0.208 ps=1.59 w=1.26 l=0.15
X83 clkb a_2432_n962# vdd vdd sky130_fd_pr__pfet_01v8 ad=0.208 pd=1.59 as=0.208 ps=1.59 w=1.26 l=0.15
X84 vdd a_2020_n482# a_2432_n962# vdd sky130_fd_pr__pfet_01v8 ad=0.208 pd=1.59 as=0.208 ps=1.59 w=1.26 l=0.15
X85 vdd a_2432_n962# clkb vdd sky130_fd_pr__pfet_01v8 ad=0.208 pd=1.59 as=0.208 ps=1.59 w=1.26 l=0.15
X86 a_2432_n962# a_2020_n482# gnd gnd sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X87 a_344_102# a_1394_n918# gnd gnd sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X88 a_2020_n482# a_344_102# vdd vdd sky130_fd_pr__pfet_01v8 ad=0.208 pd=1.59 as=0.391 ps=3.14 w=1.26 l=0.15
X89 clkb a_2432_n962# gnd gnd sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X90 gnd a_344_102# a_2020_n482# gnd sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X91 a_992_n918# a_786_n912# gnd gnd sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X92 gnd a_2432_n962# clkb gnd sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X93 clkb a_2432_n962# vdd vdd sky130_fd_pr__pfet_01v8 ad=0.391 pd=3.14 as=0.208 ps=1.59 w=1.26 l=0.15
X94 vdd a_2432_n962# clkb vdd sky130_fd_pr__pfet_01v8 ad=0.208 pd=1.59 as=0.208 ps=1.59 w=1.26 l=0.15
X95 clkb a_2432_n962# gnd gnd sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X96 a_786_n2# a_586_n2# vdd vdd sky130_fd_pr__pfet_01v8 ad=0.365 pd=3.1 as=0.365 ps=3.1 w=1.26 l=0.15
X97 clkb a_2432_n962# vdd vdd sky130_fd_pr__pfet_01v8 ad=0.208 pd=1.59 as=0.208 ps=1.59 w=1.26 l=0.15
C0 clkb vdd 7.31f
C1 a_2432_n962# clkb 2.67f
C2 a_2020_n482# vdd 2.66f
C3 a_2432_n962# vdd 7.04f
C4 clkb gnd 5.1f
C5 a_2432_n962# gnd 8.71f
C6 a_2020_n482# gnd 2.57f
C7 vdd gnd 26.1f
C8 a_344_102# gnd 2.81f
C9 a_2402_572# gnd 2.31f
C10 a_344_n986# gnd 2.43f
C11 a_3246_118# gnd 6.79f
.ends

.subckt buffer_digital i in VDD GND
Xsky130_fd_pr__pfet_01v8_FXZ64Q_0 VDD VDD a_116_148# i GND sky130_fd_pr__pfet_01v8_FXZ64Q
Xsky130_fd_pr__pfet_01v8_FXZ64Q_1 VDD VDD in a_116_148# GND sky130_fd_pr__pfet_01v8_FXZ64Q
Xsky130_fd_pr__nfet_01v8_DQBD8A_0 a_116_148# i GND GND sky130_fd_pr__nfet_01v8_DQBD8A
Xsky130_fd_pr__nfet_01v8_DQBD8A_1 in a_116_148# GND GND sky130_fd_pr__nfet_01v8_DQBD8A
.ends

.subckt sky130_fd_pr__pfet_01v8_4ZKXAA a_63_n42# a_n417_n42# a_303_n139# w_n545_n142#
+ a_255_n42# a_n465_n139# a_n129_n42# a_111_n139# a_447_n42# a_n273_n139# a_n177_73#
+ a_n321_n42# a_207_73# a_n509_n42# a_159_n42# a_15_73# a_n81_n139# a_351_n42# a_n33_n42#
+ a_n369_73# a_n225_n42# a_399_73# VSUBS
X0 a_n33_n42# a_n81_n139# a_n129_n42# w_n545_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X1 a_351_n42# a_303_n139# a_255_n42# w_n545_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X2 a_159_n42# a_111_n139# a_63_n42# w_n545_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X3 a_255_n42# a_207_73# a_159_n42# w_n545_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X4 a_447_n42# a_399_73# a_351_n42# w_n545_n142# sky130_fd_pr__pfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X5 a_n321_n42# a_n369_73# a_n417_n42# w_n545_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X6 a_n225_n42# a_n273_n139# a_n321_n42# w_n545_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X7 a_n417_n42# a_n465_n139# a_n509_n42# w_n545_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X8 a_n129_n42# a_n177_73# a_n225_n42# w_n545_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X9 a_63_n42# a_15_73# a_n33_n42# w_n545_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
.ends

.subckt sky130_fd_pr__nfet_01v8_9LGCGE a_15_n130# a_n561_n130# a_63_n42# a_n989_n42#
+ a_n177_n130# a_n417_n42# a_n465_64# a_255_n42# a_495_64# a_735_n42# a_n129_n42#
+ a_n609_n42# a_111_64# a_447_n42# a_927_n42# a_783_n130# a_n321_n42# a_399_n130#
+ a_n657_64# a_n801_n42# a_687_64# a_n945_n130# a_159_n42# a_639_n42# a_n513_n42#
+ a_n897_n42# a_591_n130# a_n81_64# a_n273_64# a_351_n42# a_207_n130# a_303_64# a_n33_n42#
+ a_831_n42# a_n369_n130# a_n753_n130# a_n849_64# a_n225_n42# a_n705_n42# a_879_64#
+ a_543_n42# VSUBS
X0 a_63_n42# a_15_n130# a_n33_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X1 a_927_n42# a_879_64# a_831_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X2 a_n33_n42# a_n81_64# a_n129_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X3 a_351_n42# a_303_64# a_255_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X4 a_159_n42# a_111_64# a_63_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X5 a_255_n42# a_207_n130# a_159_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X6 a_447_n42# a_399_n130# a_351_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X7 a_543_n42# a_495_64# a_447_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X8 a_735_n42# a_687_64# a_639_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X9 a_831_n42# a_783_n130# a_735_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X10 a_639_n42# a_591_n130# a_543_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X11 a_n321_n42# a_n369_n130# a_n417_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X12 a_n801_n42# a_n849_64# a_n897_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X13 a_n705_n42# a_n753_n130# a_n801_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X14 a_n609_n42# a_n657_64# a_n705_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X15 a_n513_n42# a_n561_n130# a_n609_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X16 a_n417_n42# a_n465_64# a_n513_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X17 a_n225_n42# a_n273_64# a_n321_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X18 a_n129_n42# a_n177_n130# a_n225_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X19 a_n897_n42# a_n945_n130# a_n989_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
.ends

.subckt sky130_fd_pr__pfet_01v8_49FP49 a_63_n42# a_n989_n42# a_n369_n139# a_n753_n139#
+ a_n417_n42# a_687_73# w_n1025_n142# a_255_n42# a_735_n42# a_n81_73# a_n273_73# a_n129_n42#
+ a_15_n139# a_n561_n139# a_303_73# a_n609_n42# a_n177_n139# a_n849_73# a_447_n42#
+ a_927_n42# a_n321_n42# a_879_73# a_n801_n42# a_159_n42# a_639_n42# a_n465_73# a_n513_n42#
+ a_n897_n42# a_783_n139# a_495_73# a_399_n139# a_351_n42# a_n33_n42# a_831_n42# a_n945_n139#
+ a_n225_n42# a_n705_n42# a_111_73# a_591_n139# a_543_n42# a_207_n139# a_n657_73#
+ VSUBS
X0 a_927_n42# a_879_73# a_831_n42# w_n1025_n142# sky130_fd_pr__pfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X1 a_n33_n42# a_n81_73# a_n129_n42# w_n1025_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X2 a_351_n42# a_303_73# a_255_n42# w_n1025_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X3 a_159_n42# a_111_73# a_63_n42# w_n1025_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X4 a_255_n42# a_207_n139# a_159_n42# w_n1025_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X5 a_447_n42# a_399_n139# a_351_n42# w_n1025_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X6 a_543_n42# a_495_73# a_447_n42# w_n1025_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X7 a_639_n42# a_591_n139# a_543_n42# w_n1025_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X8 a_735_n42# a_687_73# a_639_n42# w_n1025_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X9 a_831_n42# a_783_n139# a_735_n42# w_n1025_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X10 a_n801_n42# a_n849_73# a_n897_n42# w_n1025_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X11 a_n513_n42# a_n561_n139# a_n609_n42# w_n1025_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X12 a_n321_n42# a_n369_n139# a_n417_n42# w_n1025_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X13 a_n225_n42# a_n273_73# a_n321_n42# w_n1025_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X14 a_n897_n42# a_n945_n139# a_n989_n42# w_n1025_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X15 a_n705_n42# a_n753_n139# a_n801_n42# w_n1025_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X16 a_n609_n42# a_n657_73# a_n705_n42# w_n1025_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X17 a_n417_n42# a_n465_73# a_n513_n42# w_n1025_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X18 a_n129_n42# a_n177_n139# a_n225_n42# w_n1025_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X19 a_63_n42# a_15_n139# a_n33_n42# w_n1025_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
.ends

.subckt sky130_fd_pr__nfet_01v8_NJGC45 a_63_n42# a_15_64# a_n417_n42# a_111_n130#
+ a_n273_n130# a_255_n42# a_n129_n42# a_n369_64# a_399_64# a_447_n42# a_n81_n130#
+ a_n321_n42# a_n509_n42# a_159_n42# a_351_n42# a_n33_n42# a_303_n130# a_n225_n42#
+ a_n177_64# a_207_64# a_n465_n130# VSUBS
X0 a_63_n42# a_15_64# a_n33_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X1 a_n33_n42# a_n81_n130# a_n129_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X2 a_351_n42# a_303_n130# a_255_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X3 a_159_n42# a_111_n130# a_63_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X4 a_255_n42# a_207_64# a_159_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X5 a_447_n42# a_399_64# a_351_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X6 a_n321_n42# a_n369_64# a_n417_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X7 a_n417_n42# a_n465_n130# a_n509_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X8 a_n225_n42# a_n273_n130# a_n321_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X9 a_n129_n42# a_n177_64# a_n225_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
.ends

.subckt buffer a_1504_1398# m5_n1320_776# a_n1158_1778# a_1504_1860# a_1596_1398#
+ sky130_fd_pr__pfet_01v8_VR4B8J_1/VSUBS w_1358_2156# m4_n1330_2222#
Xsky130_fd_pr__nfet_01v8_NJGLN5_1 a_n1158_1778# sky130_fd_pr__pfet_01v8_VR4B8J_1/VSUBS
+ a_n1158_1778# a_n1158_1778# a_n1158_1778# a_n1158_1778# a_n1158_1778# a_1436_1552#
+ a_n1158_1778# a_n1158_1778# a_1436_1552# a_1436_1552# sky130_fd_pr__pfet_01v8_VR4B8J_1/VSUBS
+ sky130_fd_pr__pfet_01v8_VR4B8J_1/VSUBS a_n1158_1778# a_1436_1552# a_n1158_1778#
+ a_n1158_1778# a_n1158_1778# a_n1158_1778# a_1436_1552# sky130_fd_pr__pfet_01v8_VR4B8J_1/VSUBS
+ a_1436_1552# a_1436_1552# a_n1158_1778# sky130_fd_pr__pfet_01v8_VR4B8J_1/VSUBS sky130_fd_pr__pfet_01v8_VR4B8J_1/VSUBS
+ a_n1158_1778# a_1436_1552# a_n1158_1778# a_n1158_1778# a_n1158_1778# a_1436_1552#
+ sky130_fd_pr__pfet_01v8_VR4B8J_1/VSUBS a_n1158_1778# a_n1158_1778# sky130_fd_pr__pfet_01v8_VR4B8J_1/VSUBS
+ a_1436_1552# sky130_fd_pr__pfet_01v8_VR4B8J_1/VSUBS a_n1158_1778# sky130_fd_pr__pfet_01v8_VR4B8J_1/VSUBS
+ a_n1158_1778# a_n1158_1778# a_n1158_1778# a_n1158_1778# a_1436_1552# a_n1158_1778#
+ sky130_fd_pr__pfet_01v8_VR4B8J_1/VSUBS a_1436_1552# sky130_fd_pr__pfet_01v8_VR4B8J_1/VSUBS
+ sky130_fd_pr__pfet_01v8_VR4B8J_1/VSUBS a_1436_1552# a_1436_1552# sky130_fd_pr__pfet_01v8_VR4B8J_1/VSUBS
+ a_n1158_1778# sky130_fd_pr__pfet_01v8_VR4B8J_1/VSUBS sky130_fd_pr__nfet_01v8_NJGLN5
Xsky130_fd_pr__pfet_01v8_VR4B8J_1 a_n1158_1778# w_1358_2156# a_1436_1552# a_1436_1552#
+ w_1358_2156# a_1436_1552# a_n1158_1778# a_1436_1552# w_1358_2156# a_n1158_1778#
+ a_n1158_1778# a_n1158_1778# a_n1158_1778# a_n1158_1778# a_n1158_1778# a_n1158_1778#
+ w_1358_2156# a_1436_1552# w_1358_2156# a_n1158_1778# w_1358_2156# w_1358_2156# w_1358_2156#
+ a_n1158_1778# a_1436_1552# a_n1158_1778# a_n1158_1778# a_n1158_1778# a_n1158_1778#
+ a_1436_1552# w_1358_2156# a_n1158_1778# w_1358_2156# w_1358_2156# a_n1158_1778#
+ w_1358_2156# a_n1158_1778# w_1358_2156# a_1436_1552# a_1436_1552# a_1436_1552# a_n1158_1778#
+ a_n1158_1778# a_n1158_1778# a_1436_1552# w_1358_2156# w_1358_2156# a_n1158_1778#
+ a_n1158_1778# a_1436_1552# a_n1158_1778# a_1436_1552# a_1436_1552# a_n1158_1778#
+ a_n1158_1778# a_n1158_1778# sky130_fd_pr__pfet_01v8_VR4B8J_1/VSUBS sky130_fd_pr__pfet_01v8_VR4B8J
X0 a_1504_1398# a_1436_1552# a_1596_1398# sky130_fd_pr__pfet_01v8_VR4B8J_1/VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X1 a_1504_1860# a_1436_1552# a_1596_1398# w_1358_2156# sky130_fd_pr__pfet_01v8 ad=0.208 pd=1.59 as=0.208 ps=1.59 w=1.26 l=0.15
X2 a_1596_1398# a_1436_1552# a_1504_1398# sky130_fd_pr__pfet_01v8_VR4B8J_1/VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X3 a_1596_1398# a_1436_1552# a_1504_1860# w_1358_2156# sky130_fd_pr__pfet_01v8 ad=0.208 pd=1.59 as=0.208 ps=1.59 w=1.26 l=0.15
X4 a_1596_1398# a_1436_1552# a_1504_1860# w_1358_2156# sky130_fd_pr__pfet_01v8 ad=0.391 pd=3.14 as=0.208 ps=1.59 w=1.26 l=0.15
X5 a_1596_1398# a_1436_1552# a_1504_1860# w_1358_2156# sky130_fd_pr__pfet_01v8 ad=0.208 pd=1.59 as=0.391 ps=3.14 w=1.26 l=0.15
X6 a_1596_1398# a_1436_1552# a_1504_1398# sky130_fd_pr__pfet_01v8_VR4B8J_1/VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X7 a_1504_1860# a_1436_1552# a_1596_1398# w_1358_2156# sky130_fd_pr__pfet_01v8 ad=0.208 pd=1.59 as=0.208 ps=1.59 w=1.26 l=0.15
X8 a_1596_1398# a_1436_1552# a_1504_1398# sky130_fd_pr__pfet_01v8_VR4B8J_1/VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X9 a_1504_1398# a_1436_1552# a_1596_1398# sky130_fd_pr__pfet_01v8_VR4B8J_1/VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X10 a_1504_1860# a_1436_1552# a_1596_1398# w_1358_2156# sky130_fd_pr__pfet_01v8 ad=0.208 pd=1.59 as=0.208 ps=1.59 w=1.26 l=0.15
X11 a_1596_1398# a_1436_1552# a_1504_1860# w_1358_2156# sky130_fd_pr__pfet_01v8 ad=0.208 pd=1.59 as=0.208 ps=1.59 w=1.26 l=0.15
X12 a_1504_1398# a_1436_1552# a_1596_1398# sky130_fd_pr__pfet_01v8_VR4B8J_1/VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X13 a_1596_1398# a_1436_1552# a_1504_1398# sky130_fd_pr__pfet_01v8_VR4B8J_1/VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X14 a_1596_1398# a_1436_1552# a_1504_1860# w_1358_2156# sky130_fd_pr__pfet_01v8 ad=0.208 pd=1.59 as=0.208 ps=1.59 w=1.26 l=0.15
X15 a_1504_1860# a_1436_1552# a_1596_1398# w_1358_2156# sky130_fd_pr__pfet_01v8 ad=0.208 pd=1.59 as=0.208 ps=1.59 w=1.26 l=0.15
X16 a_1504_1860# a_1436_1552# a_1596_1398# w_1358_2156# sky130_fd_pr__pfet_01v8 ad=0.208 pd=1.59 as=0.208 ps=1.59 w=1.26 l=0.15
X17 a_1504_1398# a_1436_1552# a_1596_1398# sky130_fd_pr__pfet_01v8_VR4B8J_1/VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X18 a_1596_1398# a_1436_1552# a_1504_1398# sky130_fd_pr__pfet_01v8_VR4B8J_1/VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X19 a_1596_1398# a_1436_1552# a_1504_1860# w_1358_2156# sky130_fd_pr__pfet_01v8 ad=0.208 pd=1.59 as=0.208 ps=1.59 w=1.26 l=0.15
X20 a_1596_1398# a_1436_1552# a_1504_1860# w_1358_2156# sky130_fd_pr__pfet_01v8 ad=0.208 pd=1.59 as=0.208 ps=1.59 w=1.26 l=0.15
X21 a_1504_1398# a_1436_1552# a_1596_1398# sky130_fd_pr__pfet_01v8_VR4B8J_1/VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X22 a_1596_1398# a_1436_1552# a_1504_1398# sky130_fd_pr__pfet_01v8_VR4B8J_1/VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X23 a_1504_1860# a_1436_1552# a_1596_1398# w_1358_2156# sky130_fd_pr__pfet_01v8 ad=0.208 pd=1.59 as=0.208 ps=1.59 w=1.26 l=0.15
X24 a_1504_1398# a_1436_1552# a_1596_1398# sky130_fd_pr__pfet_01v8_VR4B8J_1/VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X25 a_1504_1398# a_1436_1552# a_1596_1398# sky130_fd_pr__pfet_01v8_VR4B8J_1/VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X26 a_1596_1398# a_1436_1552# a_1504_1860# w_1358_2156# sky130_fd_pr__pfet_01v8 ad=0.208 pd=1.59 as=0.208 ps=1.59 w=1.26 l=0.15
X27 a_1596_1398# a_1436_1552# a_1504_1398# sky130_fd_pr__pfet_01v8_VR4B8J_1/VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X28 a_1504_1398# a_1436_1552# a_1596_1398# sky130_fd_pr__pfet_01v8_VR4B8J_1/VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X29 a_1596_1398# a_1436_1552# a_1504_1860# w_1358_2156# sky130_fd_pr__pfet_01v8 ad=0.208 pd=1.59 as=0.208 ps=1.59 w=1.26 l=0.15
X30 a_1504_1398# a_1436_1552# a_1596_1398# sky130_fd_pr__pfet_01v8_VR4B8J_1/VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X31 a_1596_1398# a_1436_1552# a_1504_1860# w_1358_2156# sky130_fd_pr__pfet_01v8 ad=0.208 pd=1.59 as=0.208 ps=1.59 w=1.26 l=0.15
X32 a_1596_1398# a_1436_1552# a_1504_1398# sky130_fd_pr__pfet_01v8_VR4B8J_1/VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X33 a_1596_1398# a_1436_1552# a_1504_1398# sky130_fd_pr__pfet_01v8_VR4B8J_1/VSUBS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X34 a_1504_1860# a_1436_1552# a_1596_1398# w_1358_2156# sky130_fd_pr__pfet_01v8 ad=0.208 pd=1.59 as=0.208 ps=1.59 w=1.26 l=0.15
X35 a_1596_1398# a_1436_1552# a_1504_1398# sky130_fd_pr__pfet_01v8_VR4B8J_1/VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X36 a_1504_1398# a_1436_1552# a_1596_1398# sky130_fd_pr__pfet_01v8_VR4B8J_1/VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X37 a_1504_1860# a_1436_1552# a_1596_1398# w_1358_2156# sky130_fd_pr__pfet_01v8 ad=0.208 pd=1.59 as=0.208 ps=1.59 w=1.26 l=0.15
X38 a_1596_1398# a_1436_1552# a_1504_1860# w_1358_2156# sky130_fd_pr__pfet_01v8 ad=0.208 pd=1.59 as=0.208 ps=1.59 w=1.26 l=0.15
X39 a_1504_1398# a_1436_1552# a_1596_1398# sky130_fd_pr__pfet_01v8_VR4B8J_1/VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X40 a_1596_1398# a_1436_1552# a_1504_1398# sky130_fd_pr__pfet_01v8_VR4B8J_1/VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X41 a_1596_1398# a_1436_1552# a_1504_1398# sky130_fd_pr__pfet_01v8_VR4B8J_1/VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X42 a_1504_1860# a_1436_1552# a_1596_1398# w_1358_2156# sky130_fd_pr__pfet_01v8 ad=0.208 pd=1.59 as=0.208 ps=1.59 w=1.26 l=0.15
X43 a_1504_1398# a_1436_1552# a_1596_1398# sky130_fd_pr__pfet_01v8_VR4B8J_1/VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X44 a_1596_1398# a_1436_1552# a_1504_1860# w_1358_2156# sky130_fd_pr__pfet_01v8 ad=0.208 pd=1.59 as=0.208 ps=1.59 w=1.26 l=0.15
X45 a_1504_1860# a_1436_1552# a_1596_1398# w_1358_2156# sky130_fd_pr__pfet_01v8 ad=0.208 pd=1.59 as=0.208 ps=1.59 w=1.26 l=0.15
X46 a_1504_1398# a_1436_1552# a_1596_1398# sky130_fd_pr__pfet_01v8_VR4B8J_1/VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X47 a_1596_1398# a_1436_1552# a_1504_1860# w_1358_2156# sky130_fd_pr__pfet_01v8 ad=0.208 pd=1.59 as=0.208 ps=1.59 w=1.26 l=0.15
X48 a_1504_1860# a_1436_1552# a_1596_1398# w_1358_2156# sky130_fd_pr__pfet_01v8 ad=0.208 pd=1.59 as=0.208 ps=1.59 w=1.26 l=0.15
X49 a_1504_1860# a_1436_1552# a_1596_1398# w_1358_2156# sky130_fd_pr__pfet_01v8 ad=0.208 pd=1.59 as=0.208 ps=1.59 w=1.26 l=0.15
X50 a_1596_1398# a_1436_1552# a_1504_1398# sky130_fd_pr__pfet_01v8_VR4B8J_1/VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X51 a_1596_1398# a_1436_1552# a_1504_1398# sky130_fd_pr__pfet_01v8_VR4B8J_1/VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X52 a_1596_1398# a_1436_1552# a_1504_1860# w_1358_2156# sky130_fd_pr__pfet_01v8 ad=0.208 pd=1.59 as=0.208 ps=1.59 w=1.26 l=0.15
X53 a_1504_1860# a_1436_1552# a_1596_1398# w_1358_2156# sky130_fd_pr__pfet_01v8 ad=0.208 pd=1.59 as=0.208 ps=1.59 w=1.26 l=0.15
C0 a_1436_1552# w_1358_2156# 4.34f
C1 a_1596_1398# a_1436_1552# 2.21f
C2 a_1596_1398# a_1504_1398# 2.65f
C3 a_1596_1398# a_1504_1860# 6.79f
C4 m5_n1320_776# sky130_fd_pr__pfet_01v8_VR4B8J_1/VSUBS 2.59f
C5 a_n1158_1778# sky130_fd_pr__pfet_01v8_VR4B8J_1/VSUBS 8.21f
C6 w_1358_2156# sky130_fd_pr__pfet_01v8_VR4B8J_1/VSUBS 6.12f
C7 a_1436_1552# sky130_fd_pr__pfet_01v8_VR4B8J_1/VSUBS 9.83f
.ends

.subckt sky130_fd_pr__pfet_01v8_X4L24Q a_n33_n126# w_n353_n226# a_n317_n126# a_n177_157#
+ a_159_n126# a_111_n223# a_n273_n223# a_255_n126# a_n129_n126# a_n81_n223# a_63_n126#
+ a_n225_n126# a_15_157# a_207_157# VSUBS
X0 a_159_n126# a_111_n223# a_63_n126# w_n353_n226# sky130_fd_pr__pfet_01v8 ad=0.208 pd=1.59 as=0.208 ps=1.59 w=1.26 l=0.15
X1 a_n225_n126# a_n273_n223# a_n317_n126# w_n353_n226# sky130_fd_pr__pfet_01v8 ad=0.208 pd=1.59 as=0.391 ps=3.14 w=1.26 l=0.15
X2 a_63_n126# a_15_157# a_n33_n126# w_n353_n226# sky130_fd_pr__pfet_01v8 ad=0.208 pd=1.59 as=0.208 ps=1.59 w=1.26 l=0.15
X3 a_n129_n126# a_n177_157# a_n225_n126# w_n353_n226# sky130_fd_pr__pfet_01v8 ad=0.208 pd=1.59 as=0.208 ps=1.59 w=1.26 l=0.15
X4 a_n33_n126# a_n81_n223# a_n129_n126# w_n353_n226# sky130_fd_pr__pfet_01v8 ad=0.208 pd=1.59 as=0.208 ps=1.59 w=1.26 l=0.15
X5 a_255_n126# a_207_157# a_159_n126# w_n353_n226# sky130_fd_pr__pfet_01v8 ad=0.391 pd=3.14 as=0.208 ps=1.59 w=1.26 l=0.15
.ends

.subckt sky130_fd_pr__nfet_01v8_XJUN3E a_63_n42# a_15_64# a_111_n130# a_n273_n130#
+ a_255_n42# a_n129_n42# a_n317_n42# a_n81_n130# a_159_n42# a_n33_n42# a_n225_n42#
+ a_n177_64# a_207_64# VSUBS
X0 a_63_n42# a_15_64# a_n33_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X1 a_n33_n42# a_n81_n130# a_n129_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X2 a_159_n42# a_111_n130# a_63_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X3 a_255_n42# a_207_64# a_159_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X4 a_n225_n42# a_n273_n130# a_n317_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X5 a_n129_n42# a_n177_64# a_n225_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
.ends

.subckt and_gate a_514_134# w_n260_286# sky130_fd_pr__pfet_01v8_X4L24Q_0/VSUBS a_n162_206#
+ m1_748_n50#
Xsky130_fd_pr__pfet_01v8_X4L24Q_0 w_n260_286# w_n260_286# m1_748_n50# a_n78_396# w_n260_286#
+ a_n78_396# a_n78_396# m1_748_n50# m1_748_n50# a_n78_396# m1_748_n50# w_n260_286#
+ a_n78_396# a_n78_396# sky130_fd_pr__pfet_01v8_X4L24Q_0/VSUBS sky130_fd_pr__pfet_01v8_X4L24Q
Xsky130_fd_pr__nfet_01v8_XJUN3E_0 m1_748_n50# a_n78_396# a_n78_396# a_n78_396# m1_748_n50#
+ m1_748_n50# m1_748_n50# a_n78_396# sky130_fd_pr__pfet_01v8_X4L24Q_0/VSUBS sky130_fd_pr__pfet_01v8_X4L24Q_0/VSUBS
+ sky130_fd_pr__pfet_01v8_X4L24Q_0/VSUBS a_n78_396# a_n78_396# sky130_fd_pr__pfet_01v8_X4L24Q_0/VSUBS
+ sky130_fd_pr__nfet_01v8_XJUN3E
X0 a_n78_396# a_n162_206# w_n260_286# w_n260_286# sky130_fd_pr__pfet_01v8 ad=0.208 pd=1.59 as=0.208 ps=1.59 w=1.26 l=0.15
X1 sky130_fd_pr__pfet_01v8_X4L24Q_0/VSUBS a_n162_206# a_n78_n64# sky130_fd_pr__pfet_01v8_X4L24Q_0/VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X2 w_n260_286# a_n162_206# a_n78_396# w_n260_286# sky130_fd_pr__pfet_01v8 ad=0.208 pd=1.59 as=0.208 ps=1.59 w=1.26 l=0.15
X3 w_n260_286# a_n162_206# a_n78_396# w_n260_286# sky130_fd_pr__pfet_01v8 ad=0.208 pd=1.59 as=0.208 ps=1.59 w=1.26 l=0.15
X4 a_n78_396# a_n162_206# w_n260_286# w_n260_286# sky130_fd_pr__pfet_01v8 ad=0.195 pd=1.57 as=0.208 ps=1.59 w=1.26 l=0.15
X5 a_n78_396# a_514_134# a_n78_n64# sky130_fd_pr__pfet_01v8_X4L24Q_0/VSUBS sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0651 ps=0.73 w=0.42 l=0.15
X6 a_n78_n64# a_n162_206# sky130_fd_pr__pfet_01v8_X4L24Q_0/VSUBS sky130_fd_pr__pfet_01v8_X4L24Q_0/VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X7 w_n260_286# a_514_134# a_n78_396# w_n260_286# sky130_fd_pr__pfet_01v8 ad=0.365 pd=3.1 as=0.195 ps=1.57 w=1.26 l=0.15
X8 a_n78_396# a_n162_206# w_n260_286# w_n260_286# sky130_fd_pr__pfet_01v8 ad=0.208 pd=1.59 as=0.208 ps=1.59 w=1.26 l=0.15
X9 sky130_fd_pr__pfet_01v8_X4L24Q_0/VSUBS a_n162_206# a_n78_n64# sky130_fd_pr__pfet_01v8_X4L24Q_0/VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X10 w_n260_286# a_n162_206# a_n78_396# w_n260_286# sky130_fd_pr__pfet_01v8 ad=0.208 pd=1.59 as=0.391 ps=3.14 w=1.26 l=0.15
X11 sky130_fd_pr__pfet_01v8_X4L24Q_0/VSUBS a_n162_206# a_n78_n64# sky130_fd_pr__pfet_01v8_X4L24Q_0/VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X12 a_n78_n64# a_n162_206# sky130_fd_pr__pfet_01v8_X4L24Q_0/VSUBS sky130_fd_pr__pfet_01v8_X4L24Q_0/VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X13 a_n78_n64# a_n162_206# sky130_fd_pr__pfet_01v8_X4L24Q_0/VSUBS sky130_fd_pr__pfet_01v8_X4L24Q_0/VSUBS sky130_fd_pr__nfet_01v8 ad=0.0651 pd=0.73 as=0.0693 ps=0.75 w=0.42 l=0.15
C0 a_n78_396# w_n260_286# 3.02f
C1 a_n78_396# sky130_fd_pr__pfet_01v8_X4L24Q_0/VSUBS 2.46f
C2 w_n260_286# sky130_fd_pr__pfet_01v8_X4L24Q_0/VSUBS 6.96f
.ends

.subckt buffer_and_gate in1 clk out gnd vdd
Xbuffer_0 gnd gnd clk vdd m1_5444_838# gnd vdd vdd buffer
Xand_gate_0 m1_5444_838# vdd gnd in1 out and_gate
C0 in1 gnd 2.62f
C1 and_gate_0/a_n78_396# gnd 2.34f
C2 clk gnd 8.8f
C3 m1_5444_838# gnd 2.35f
C4 vdd gnd 18.3f
C5 buffer_0/a_1436_1552# gnd 11.5f
.ends

.subckt capacito7 a_2858_n174# sky130_fd_pr__pfet_01v8_4ZKXAA_0/w_n545_n142# buffer_digital_0/i
+ a_5270_n124# m3_7758_166# buffer_and_gate_0/clk sky130_fd_pr__pfet_01v8_49FP49_0/w_n1025_n142#
+ m1_6370_n278# buffer_digital_0/VDD m1_602_n334# VSUBS
Xbuffer_digital_0 buffer_digital_0/i buffer_digital_0/in buffer_digital_0/VDD VSUBS
+ buffer_digital
Xsky130_fd_pr__pfet_01v8_4ZKXAA_0 m1_6370_n278# m1_6370_n278# VSUBS sky130_fd_pr__pfet_01v8_4ZKXAA_0/w_n545_n142#
+ m1_6370_n278# VSUBS m1_6370_n278# VSUBS m1_6370_n278# VSUBS VSUBS m1_6370_n278#
+ VSUBS m1_6370_n278# m1_6370_n278# VSUBS VSUBS m1_6370_n278# m1_6370_n278# VSUBS
+ m1_6370_n278# VSUBS VSUBS sky130_fd_pr__pfet_01v8_4ZKXAA
Xsky130_fd_pr__nfet_01v8_9LGCGE_0 a_2858_n174# a_2858_n174# VSUBS VSUBS a_2858_n174#
+ VSUBS a_2858_n174# VSUBS a_2858_n174# VSUBS VSUBS VSUBS a_2858_n174# VSUBS VSUBS
+ a_2858_n174# VSUBS a_2858_n174# a_2858_n174# VSUBS a_2858_n174# a_2858_n174# VSUBS
+ VSUBS VSUBS VSUBS a_2858_n174# a_2858_n174# a_2858_n174# VSUBS a_2858_n174# a_2858_n174#
+ VSUBS VSUBS a_2858_n174# a_2858_n174# a_2858_n174# VSUBS VSUBS a_2858_n174# VSUBS
+ VSUBS sky130_fd_pr__nfet_01v8_9LGCGE
Xsky130_fd_pr__pfet_01v8_49FP49_0 m1_602_n334# m1_602_n334# VSUBS VSUBS m1_602_n334#
+ VSUBS sky130_fd_pr__pfet_01v8_49FP49_0/w_n1025_n142# m1_602_n334# m1_602_n334# VSUBS
+ VSUBS m1_602_n334# VSUBS VSUBS VSUBS m1_602_n334# VSUBS VSUBS m1_602_n334# m1_602_n334#
+ m1_602_n334# VSUBS m1_602_n334# m1_602_n334# m1_602_n334# VSUBS m1_602_n334# m1_602_n334#
+ VSUBS VSUBS VSUBS m1_602_n334# m1_602_n334# m1_602_n334# VSUBS m1_602_n334# m1_602_n334#
+ VSUBS VSUBS m1_602_n334# VSUBS VSUBS VSUBS sky130_fd_pr__pfet_01v8_49FP49
Xsky130_fd_pr__nfet_01v8_NJGC45_0 VSUBS a_5270_n124# VSUBS a_5270_n124# a_5270_n124#
+ VSUBS VSUBS a_5270_n124# a_5270_n124# VSUBS a_5270_n124# VSUBS VSUBS VSUBS VSUBS
+ VSUBS a_5270_n124# VSUBS a_5270_n124# a_5270_n124# a_5270_n124# VSUBS sky130_fd_pr__nfet_01v8_NJGC45
Xbuffer_and_gate_0 buffer_digital_0/in buffer_and_gate_0/clk buffer_and_gate_0/out
+ VSUBS buffer_digital_0/VDD buffer_and_gate
X0 buffer_and_gate_0/out m3_7758_166# sky130_fd_pr__cap_mim_m3_1 l=7.99 w=7.97
C0 buffer_digital_0/i buffer_digital_0/in 2.94f
C1 m3_7758_166# VSUBS 2.5f
C2 buffer_and_gate_0/and_gate_0/a_n78_396# VSUBS 2.47f
C3 buffer_and_gate_0/clk VSUBS 8.92f
C4 buffer_digital_0/VDD VSUBS 18f
C5 buffer_and_gate_0/buffer_0/a_1436_1552# VSUBS 10.2f
C6 a_5270_n124# VSUBS 3.42f
C7 m1_602_n334# VSUBS 2.78f
C8 a_2858_n174# VSUBS 6.7f
C9 buffer_digital_0/in VSUBS 2.68f
.ends

.subckt capacitor_8 capacitor_7_0/a_5270_n124# capacitor_7_0/m3_7758_166# capacitor_7_0/buffer_and_gate_0/clk
+ capacitor_7_0/buffer_digital_0/VDD capacitor_7_0/a_2858_n174# w_7118_n356# w_1380_n364#
+ VSUBS capacitor_7_0/buffer_digital_0/i
Xcapacitor_7_0 capacitor_7_0/a_2858_n174# w_7118_n356# capacitor_7_0/buffer_digital_0/i
+ capacitor_7_0/a_5270_n124# capacitor_7_0/m3_7758_166# capacitor_7_0/buffer_and_gate_0/clk
+ w_1380_n364# w_7118_n356# capacitor_7_0/buffer_digital_0/VDD w_1380_n364# VSUBS
+ capacito7
C0 capacitor_7_0/m3_7758_166# VSUBS 2.32f
C1 capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# VSUBS 2.34f
C2 capacitor_7_0/buffer_and_gate_0/clk VSUBS 8.2f
C3 capacitor_7_0/buffer_digital_0/VDD VSUBS 18.2f
C4 capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# VSUBS 9.98f
C5 capacitor_7_0/a_5270_n124# VSUBS 2.36f
C6 w_1380_n364# VSUBS 3.54f
C7 capacitor_7_0/a_2858_n174# VSUBS 4.67f
C8 capacitor_7_0/buffer_digital_0/in VSUBS 2.61f
.ends

.subckt capacitors_1 clk1 capacitor_8_0/capacitor_7_0/a_2858_n174# capacitor_8_0/capacitor_7_0/a_5270_n124#
+ capacitor_8_0/capacitor_7_0/buffer_and_gate_0/clk capacitor_8_0/capacitor_7_0/buffer_digital_0/VDD
+ m1_7096_n308# capacitor_8_0/w_1380_n364# in1 VSUBS
Xcapacitor_8_0 capacitor_8_0/capacitor_7_0/a_5270_n124# clk1 capacitor_8_0/capacitor_7_0/buffer_and_gate_0/clk
+ capacitor_8_0/capacitor_7_0/buffer_digital_0/VDD capacitor_8_0/capacitor_7_0/a_2858_n174#
+ m1_7096_n308# capacitor_8_0/w_1380_n364# VSUBS in1 capacitor_8
C0 clk1 VSUBS 2.38f
C1 capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# VSUBS 2.34f
C2 capacitor_8_0/capacitor_7_0/buffer_and_gate_0/clk VSUBS 9.49f
C3 capacitor_8_0/capacitor_7_0/buffer_digital_0/VDD VSUBS 22.9f
C4 capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# VSUBS 9.98f
C5 capacitor_8_0/capacitor_7_0/a_5270_n124# VSUBS 2.36f
C6 capacitor_8_0/w_1380_n364# VSUBS 3.27f
C7 capacitor_8_0/capacitor_7_0/a_2858_n174# VSUBS 4.67f
C8 capacitor_8_0/capacitor_7_0/buffer_digital_0/in VSUBS 2.61f
.ends

.subckt sky130_fd_pr__pfet_01v8_4RPJ49 a_2031_73# a_1887_n42# a_3615_n42# a_3183_73#
+ a_n3729_73# a_n2529_n42# a_1503_n42# a_63_n42# a_n753_n139# a_n3393_n42# a_n369_n139#
+ a_n1425_73# a_n1281_n42# a_n2961_73# a_687_73# a_n2577_73# a_n417_n42# a_2367_n42#
+ a_n1761_n42# a_n3009_n42# a_n2673_n139# a_2847_n42# a_n2289_n139# a_n3633_n139#
+ a_2607_73# a_n3249_n139# a_n1713_n139# a_3759_73# a_n1329_n139# a_255_n42# a_1455_73#
+ a_n2241_n42# a_2991_73# a_3471_n139# a_735_n42# a_1551_n139# a_3087_n139# a_1599_n42#
+ a_3327_n42# a_1167_n139# a_n2721_n42# a_n81_73# a_2511_n139# a_1215_n42# a_n273_73#
+ a_2127_n139# a_n993_n42# a_3807_n42# a_15_n139# a_303_73# a_n3585_n42# a_n129_n42#
+ a_2079_n42# a_n561_n139# a_n3345_73# a_n3201_n42# a_n1473_n42# a_n177_n139# a_n1041_73#
+ a_n609_n42# a_2559_n42# a_n2193_73# a_n1953_n42# a_n849_73# w_n3905_n142# a_n2481_n139#
+ a_n2097_n139# a_n3441_n139# a_1791_n42# a_n1521_n139# a_n3057_n139# a_2223_73# a_447_n42#
+ a_3039_n42# a_n1137_n139# a_3375_73# a_n2433_n42# a_927_n42# a_1071_73# a_n1617_73#
+ a_n2913_n42# a_3519_n42# a_975_n139# a_879_73# a_n2769_73# a_n321_n42# a_1407_n42#
+ a_n3297_n42# a_2271_n42# a_n1185_n42# a_n801_n42# a_n3777_n42# a_2751_n42# a_n1665_n42#
+ a_1647_73# a_2799_73# a_3231_n42# a_159_n42# a_n2145_n42# a_n465_73# a_1983_n42#
+ a_3711_n42# a_639_n42# a_n2625_n42# a_1119_n42# a_n3537_73# a_n897_n42# a_n513_n42#
+ a_n1233_73# a_n3489_n42# a_2463_n42# a_783_n139# a_495_73# a_399_n139# a_n2385_73#
+ a_2895_n139# a_n3105_n42# a_n1377_n42# a_2943_n42# a_1935_n139# a_n1857_n42# a_351_n42#
+ a_2415_73# a_n33_n42# a_3567_73# a_831_n42# a_1695_n42# a_3423_n42# a_1263_73# a_n945_n139#
+ a_n2337_n42# a_1311_n42# a_n1809_73# a_n2817_n42# a_n3681_n42# a_n225_n42# a_2175_n42#
+ a_n2865_n139# a_n1089_n42# a_n3825_n139# a_111_73# a_n2001_73# a_n3869_n42# a_n705_n42#
+ a_2655_n42# a_n1905_n139# a_n3153_73# a_591_n139# a_1839_73# a_n1569_n42# a_3663_n139#
+ a_1743_n139# a_3279_n139# a_543_n42# a_207_n139# a_n657_73# a_1359_n139# a_2703_n139#
+ a_3135_n42# VSUBS a_2319_n139# a_n2049_n42# a_1023_n42#
X0 a_n2241_n42# a_n2289_n139# a_n2337_n42# w_n3905_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X1 a_n2913_n42# a_n2961_73# a_n3009_n42# w_n3905_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X2 a_n2721_n42# a_n2769_73# a_n2817_n42# w_n3905_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X3 a_n2625_n42# a_n2673_n139# a_n2721_n42# w_n3905_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X4 a_n2433_n42# a_n2481_n139# a_n2529_n42# w_n3905_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X5 a_n2337_n42# a_n2385_73# a_n2433_n42# w_n3905_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X6 a_n2145_n42# a_n2193_73# a_n2241_n42# w_n3905_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X7 a_n2049_n42# a_n2097_n139# a_n2145_n42# w_n3905_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X8 a_n2817_n42# a_n2865_n139# a_n2913_n42# w_n3905_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X9 a_n2529_n42# a_n2577_73# a_n2625_n42# w_n3905_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X10 a_2079_n42# a_2031_73# a_1983_n42# w_n3905_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X11 a_2175_n42# a_2127_n139# a_2079_n42# w_n3905_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X12 a_2271_n42# a_2223_73# a_2175_n42# w_n3905_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X13 a_2367_n42# a_2319_n139# a_2271_n42# w_n3905_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X14 a_2463_n42# a_2415_73# a_2367_n42# w_n3905_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X15 a_2655_n42# a_2607_73# a_2559_n42# w_n3905_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X16 a_2751_n42# a_2703_n139# a_2655_n42# w_n3905_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X17 a_2943_n42# a_2895_n139# a_2847_n42# w_n3905_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X18 a_2559_n42# a_2511_n139# a_2463_n42# w_n3905_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X19 a_2847_n42# a_2799_73# a_2751_n42# w_n3905_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X20 a_927_n42# a_879_73# a_831_n42# w_n3905_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X21 a_1023_n42# a_975_n139# a_927_n42# w_n3905_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X22 a_n1953_n42# a_n2001_73# a_n2049_n42# w_n3905_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X23 a_n1761_n42# a_n1809_73# a_n1857_n42# w_n3905_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X24 a_n1665_n42# a_n1713_n139# a_n1761_n42# w_n3905_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X25 a_n1857_n42# a_n1905_n139# a_n1953_n42# w_n3905_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X26 a_n1569_n42# a_n1617_73# a_n1665_n42# w_n3905_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X27 a_1119_n42# a_1071_73# a_1023_n42# w_n3905_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X28 a_1215_n42# a_1167_n139# a_1119_n42# w_n3905_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X29 a_1311_n42# a_1263_73# a_1215_n42# w_n3905_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X30 a_1407_n42# a_1359_n139# a_1311_n42# w_n3905_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X31 a_1503_n42# a_1455_73# a_1407_n42# w_n3905_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X32 a_1695_n42# a_1647_73# a_1599_n42# w_n3905_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X33 a_1791_n42# a_1743_n139# a_1695_n42# w_n3905_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X34 a_1599_n42# a_1551_n139# a_1503_n42# w_n3905_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X35 a_1887_n42# a_1839_73# a_1791_n42# w_n3905_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X36 a_1983_n42# a_1935_n139# a_1887_n42# w_n3905_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X37 a_n33_n42# a_n81_73# a_n129_n42# w_n3905_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X38 a_351_n42# a_303_73# a_255_n42# w_n3905_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X39 a_159_n42# a_111_73# a_63_n42# w_n3905_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X40 a_255_n42# a_207_n139# a_159_n42# w_n3905_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X41 a_447_n42# a_399_n139# a_351_n42# w_n3905_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X42 a_543_n42# a_495_73# a_447_n42# w_n3905_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X43 a_639_n42# a_591_n139# a_543_n42# w_n3905_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X44 a_735_n42# a_687_73# a_639_n42# w_n3905_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X45 a_831_n42# a_783_n139# a_735_n42# w_n3905_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X46 a_n1473_n42# a_n1521_n139# a_n1569_n42# w_n3905_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X47 a_n1377_n42# a_n1425_73# a_n1473_n42# w_n3905_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X48 a_n1281_n42# a_n1329_n139# a_n1377_n42# w_n3905_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X49 a_n1185_n42# a_n1233_73# a_n1281_n42# w_n3905_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X50 a_n1089_n42# a_n1137_n139# a_n1185_n42# w_n3905_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X51 a_n993_n42# a_n1041_73# a_n1089_n42# w_n3905_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X52 a_n801_n42# a_n849_73# a_n897_n42# w_n3905_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X53 a_n513_n42# a_n561_n139# a_n609_n42# w_n3905_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X54 a_n321_n42# a_n369_n139# a_n417_n42# w_n3905_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X55 a_n225_n42# a_n273_73# a_n321_n42# w_n3905_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X56 a_n897_n42# a_n945_n139# a_n993_n42# w_n3905_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X57 a_n705_n42# a_n753_n139# a_n801_n42# w_n3905_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X58 a_n609_n42# a_n657_73# a_n705_n42# w_n3905_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X59 a_n417_n42# a_n465_73# a_n513_n42# w_n3905_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X60 a_n129_n42# a_n177_n139# a_n225_n42# w_n3905_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X61 a_3327_n42# a_3279_n139# a_3231_n42# w_n3905_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X62 a_3423_n42# a_3375_73# a_3327_n42# w_n3905_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X63 a_3615_n42# a_3567_73# a_3519_n42# w_n3905_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X64 a_3711_n42# a_3663_n139# a_3615_n42# w_n3905_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X65 a_3519_n42# a_3471_n139# a_3423_n42# w_n3905_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X66 a_3807_n42# a_3759_73# a_3711_n42# w_n3905_n142# sky130_fd_pr__pfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X67 a_n3201_n42# a_n3249_n139# a_n3297_n42# w_n3905_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X68 a_63_n42# a_15_n139# a_n33_n42# w_n3905_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X69 a_n3681_n42# a_n3729_73# a_n3777_n42# w_n3905_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X70 a_n3585_n42# a_n3633_n139# a_n3681_n42# w_n3905_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X71 a_n3393_n42# a_n3441_n139# a_n3489_n42# w_n3905_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X72 a_n3297_n42# a_n3345_73# a_n3393_n42# w_n3905_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X73 a_n3105_n42# a_n3153_73# a_n3201_n42# w_n3905_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X74 a_n3009_n42# a_n3057_n139# a_n3105_n42# w_n3905_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X75 a_3231_n42# a_3183_73# a_3135_n42# w_n3905_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X76 a_n3777_n42# a_n3825_n139# a_n3869_n42# w_n3905_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X77 a_n3489_n42# a_n3537_73# a_n3585_n42# w_n3905_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X78 a_3039_n42# a_2991_73# a_2943_n42# w_n3905_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X79 a_3135_n42# a_3087_n139# a_3039_n42# w_n3905_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
C0 w_n3905_n142# VSUBS 6.63f
.ends

.subckt sky130_fd_pr__pfet_01v8_E9H44Q a_15_n42# a_n15_n68# w_n109_n104# a_n73_n42#
+ VSUBS
X0 a_15_n42# a_n15_n68# a_n73_n42# w_n109_n104# sky130_fd_pr__pfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
.ends

.subckt sky130_fd_pr__pfet_01v8_9AYYDL a_n158_n300# w_n194_n362# a_100_n300# a_n100_n326#
+ VSUBS
X0 a_100_n300# a_n100_n326# a_n158_n300# w_n194_n362# sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.87 ps=6.58 w=3 l=1
.ends

.subckt pmos_cp1 a_168_22# m1_532_58# w_n14_n142# a_424_18# m1_14_56# VSUBS
Xsky130_fd_pr__pfet_01v8_E9H44Q_0 w_n14_n142# a_168_22# w_n14_n142# a_424_18# VSUBS
+ sky130_fd_pr__pfet_01v8_E9H44Q
Xsky130_fd_pr__pfet_01v8_E9H44Q_1 a_168_22# a_424_18# w_n14_n142# w_n14_n142# VSUBS
+ sky130_fd_pr__pfet_01v8_E9H44Q
Xsky130_fd_pr__pfet_01v8_9AYYDL_0 m1_14_56# w_n14_n142# w_n14_n142# a_168_22# VSUBS
+ sky130_fd_pr__pfet_01v8_9AYYDL
Xsky130_fd_pr__pfet_01v8_9AYYDL_1 w_n14_n142# w_n14_n142# m1_532_58# a_424_18# VSUBS
+ sky130_fd_pr__pfet_01v8_9AYYDL
C0 w_n14_n142# VSUBS 2.47f
.ends

.subckt sky130_fd_pr__nfet_01v8_NJGC8F a_15_n130# a_1887_n42# a_3615_n42# a_1647_64#
+ a_n561_n130# a_n2529_n42# a_1503_n42# a_2799_64# a_63_n42# a_n177_n130# a_n3393_n42#
+ a_n1281_n42# a_n465_64# a_n417_n42# a_2367_n42# a_n1761_n42# a_n2481_n130# a_n3009_n42#
+ a_n2097_n130# a_n3441_n130# a_2847_n42# a_n1521_n130# a_n3057_n130# a_n3537_64#
+ a_n1137_n130# a_255_n42# a_n1233_64# a_495_64# a_n2241_n42# a_n2385_64# a_975_n130#
+ a_735_n42# a_1599_n42# a_3327_n42# a_n2721_n42# a_1215_n42# a_2415_64# a_n993_n42#
+ a_3807_n42# a_3567_64# a_n3585_n42# a_n129_n42# a_2079_n42# a_1263_64# a_n3201_n42#
+ a_n1473_n42# a_n1809_64# a_n609_n42# a_2559_n42# a_n1953_n42# a_111_64# a_n2001_64#
+ a_1791_n42# a_447_n42# a_n3153_64# a_3039_n42# a_n2433_n42# a_1839_64# a_927_n42#
+ a_n2913_n42# a_3519_n42# a_783_n130# a_399_n130# a_2895_n130# a_n321_n42# a_1407_n42#
+ a_n3297_n42# a_2271_n42# a_n657_64# a_n1185_n42# a_1935_n130# a_n801_n42# a_2031_64#
+ a_n3777_n42# a_2751_n42# a_3183_64# a_n1665_n42# a_n3729_64# a_n1425_64# a_687_64#
+ a_n2961_64# a_n945_n130# a_n2577_64# a_3231_n42# a_159_n42# a_n2145_n42# a_1983_n42#
+ a_3711_n42# a_2607_64# a_639_n42# a_n2625_n42# a_3759_64# a_n2865_n130# a_1119_n42#
+ a_n3825_n130# a_1455_64# a_n1905_n130# a_2991_64# a_n897_n42# a_591_n130# a_n513_n42#
+ a_n3489_n42# a_2463_n42# a_n3105_n42# a_n1377_n42# a_n81_64# a_n273_64# a_3663_n130#
+ a_3279_n130# a_2943_n42# a_1743_n130# a_207_n130# a_2703_n130# a_1359_n130# a_n1857_n42#
+ a_2319_n130# a_351_n42# a_303_64# a_n3345_64# a_n33_n42# a_831_n42# a_n1041_64#
+ a_1695_n42# a_3423_n42# a_n753_n130# a_n369_n130# a_n2193_64# a_n2337_n42# a_1311_n42#
+ a_n849_64# a_n2817_n42# a_n3681_n42# a_n225_n42# a_2223_64# a_n2673_n130# a_2175_n42#
+ a_3375_64# a_n2289_n130# a_n3633_n130# a_n1089_n42# a_n3249_n130# a_n1713_n130#
+ a_n3869_n42# a_n705_n42# a_2655_n42# a_1071_64# a_n1329_n130# a_n1617_64# a_n1569_n42#
+ a_879_64# a_n2769_64# a_3471_n130# a_3087_n130# a_1551_n130# a_2511_n130# a_543_n42#
+ a_1167_n130# a_3135_n42# a_2127_n130# VSUBS a_n2049_n42# a_1023_n42#
X0 a_n3201_n42# a_n3249_n130# a_n3297_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X1 a_63_n42# a_15_n130# a_n33_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X2 a_n3681_n42# a_n3729_64# a_n3777_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X3 a_n3585_n42# a_n3633_n130# a_n3681_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X4 a_n3393_n42# a_n3441_n130# a_n3489_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X5 a_n3297_n42# a_n3345_64# a_n3393_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X6 a_n3105_n42# a_n3153_64# a_n3201_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X7 a_n3009_n42# a_n3057_n130# a_n3105_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X8 a_n3777_n42# a_n3825_n130# a_n3869_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X9 a_n3489_n42# a_n3537_64# a_n3585_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X10 a_3135_n42# a_3087_n130# a_3039_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X11 a_3231_n42# a_3183_64# a_3135_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X12 a_3039_n42# a_2991_64# a_2943_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X13 a_n2241_n42# a_n2289_n130# a_n2337_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X14 a_n2913_n42# a_n2961_64# a_n3009_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X15 a_n2721_n42# a_n2769_64# a_n2817_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X16 a_n2625_n42# a_n2673_n130# a_n2721_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X17 a_n2433_n42# a_n2481_n130# a_n2529_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X18 a_n2337_n42# a_n2385_64# a_n2433_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X19 a_n2145_n42# a_n2193_64# a_n2241_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X20 a_n2049_n42# a_n2097_n130# a_n2145_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X21 a_n2817_n42# a_n2865_n130# a_n2913_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X22 a_n2529_n42# a_n2577_64# a_n2625_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X23 a_2175_n42# a_2127_n130# a_2079_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X24 a_2271_n42# a_2223_64# a_2175_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X25 a_2463_n42# a_2415_64# a_2367_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X26 a_2751_n42# a_2703_n130# a_2655_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X27 a_2079_n42# a_2031_64# a_1983_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X28 a_2367_n42# a_2319_n130# a_2271_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X29 a_2559_n42# a_2511_n130# a_2463_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X30 a_2655_n42# a_2607_64# a_2559_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X31 a_2847_n42# a_2799_64# a_2751_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X32 a_2943_n42# a_2895_n130# a_2847_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X33 a_927_n42# a_879_64# a_831_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X34 a_1023_n42# a_975_n130# a_927_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X35 a_n1953_n42# a_n2001_64# a_n2049_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X36 a_n1761_n42# a_n1809_64# a_n1857_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X37 a_n1665_n42# a_n1713_n130# a_n1761_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X38 a_n1857_n42# a_n1905_n130# a_n1953_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X39 a_n1569_n42# a_n1617_64# a_n1665_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X40 a_1215_n42# a_1167_n130# a_1119_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X41 a_1311_n42# a_1263_64# a_1215_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X42 a_1503_n42# a_1455_64# a_1407_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X43 a_1791_n42# a_1743_n130# a_1695_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X44 a_1119_n42# a_1071_64# a_1023_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X45 a_1407_n42# a_1359_n130# a_1311_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X46 a_1599_n42# a_1551_n130# a_1503_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X47 a_1695_n42# a_1647_64# a_1599_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X48 a_1887_n42# a_1839_64# a_1791_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X49 a_1983_n42# a_1935_n130# a_1887_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X50 a_n33_n42# a_n81_64# a_n129_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X51 a_351_n42# a_303_64# a_255_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X52 a_159_n42# a_111_64# a_63_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X53 a_255_n42# a_207_n130# a_159_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X54 a_447_n42# a_399_n130# a_351_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X55 a_543_n42# a_495_64# a_447_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X56 a_735_n42# a_687_64# a_639_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X57 a_831_n42# a_783_n130# a_735_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X58 a_639_n42# a_591_n130# a_543_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X59 a_n1473_n42# a_n1521_n130# a_n1569_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X60 a_n1281_n42# a_n1329_n130# a_n1377_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X61 a_n1185_n42# a_n1233_64# a_n1281_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X62 a_n993_n42# a_n1041_64# a_n1089_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X63 a_n1377_n42# a_n1425_64# a_n1473_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X64 a_n1089_n42# a_n1137_n130# a_n1185_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X65 a_n321_n42# a_n369_n130# a_n417_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X66 a_n801_n42# a_n849_64# a_n897_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X67 a_n705_n42# a_n753_n130# a_n801_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X68 a_n609_n42# a_n657_64# a_n705_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X69 a_n513_n42# a_n561_n130# a_n609_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X70 a_n417_n42# a_n465_64# a_n513_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X71 a_n225_n42# a_n273_64# a_n321_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X72 a_n129_n42# a_n177_n130# a_n225_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X73 a_n897_n42# a_n945_n130# a_n993_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X74 a_3327_n42# a_3279_n130# a_3231_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X75 a_3423_n42# a_3375_64# a_3327_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X76 a_3615_n42# a_3567_64# a_3519_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X77 a_3711_n42# a_3663_n130# a_3615_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X78 a_3519_n42# a_3471_n130# a_3423_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X79 a_3807_n42# a_3759_64# a_3711_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
.ends

.subckt charge_pump1 clk_in input1 input2 in1 in2 in6 in7 g1 g2 clk clkb m1_12464_n576#
+ a_3340_18086# in4 in3 in5 in8 vin vdd gnd
Xsky130_fd_pr__cap_mim_m3_1_MH6KF8_4 g1 clk gnd sky130_fd_pr__cap_mim_m3_1_MH6KF8
Xsky130_fd_pr__cap_mim_m3_1_MH6KF8_5 g2 clkb gnd sky130_fd_pr__cap_mim_m3_1_MH6KF8
Xnmos_dnw3_0 vin input1 input2 g1 g2 vin gnd nmos_dnw3
Xclock_0 clk_in vdd gnd clk clkb clock
Xcapacitor_8_0 vdd input1 clk vdd vdd vdd vdd gnd in8 capacitor_8
Xcapacitor_8_1 vdd input2 clkb vdd vdd vdd vdd gnd in8 capacitor_8
Xcapacitors_1_0 input1 vdd vdd clk vdd vdd vdd in1 gnd capacitors_1
Xcapacitors_1_1 input2 vdd vdd clkb vdd vdd vdd in1 gnd capacitors_1
Xcapacitors_1_2 input1 vdd vdd clk vdd vdd vdd in2 gnd capacitors_1
Xsky130_fd_pr__pfet_01v8_4RPJ49_0 gnd vdd vdd gnd gnd vdd vdd vdd gnd vdd gnd gnd
+ vdd gnd gnd gnd vdd vdd vdd vdd gnd vdd gnd gnd gnd gnd gnd gnd gnd vdd gnd vdd
+ gnd gnd vdd gnd gnd vdd vdd gnd vdd gnd gnd vdd gnd gnd vdd vdd gnd gnd vdd vdd
+ vdd gnd gnd vdd vdd gnd gnd vdd vdd gnd vdd gnd vdd gnd gnd gnd vdd gnd gnd gnd
+ vdd vdd gnd gnd vdd vdd gnd gnd vdd vdd gnd gnd gnd vdd vdd vdd vdd vdd vdd vdd
+ vdd vdd gnd gnd vdd vdd vdd gnd vdd vdd vdd vdd vdd gnd vdd vdd gnd vdd vdd gnd
+ gnd gnd gnd gnd vdd vdd vdd gnd vdd vdd gnd vdd gnd vdd vdd vdd gnd gnd vdd vdd
+ gnd vdd vdd vdd vdd gnd vdd gnd gnd gnd vdd vdd vdd gnd gnd gnd gnd vdd gnd gnd
+ gnd vdd gnd gnd gnd gnd vdd gnd gnd vdd vdd sky130_fd_pr__pfet_01v8_4RPJ49
Xcapacitors_1_3 input1 vdd vdd clk vdd vdd vdd in3 gnd capacitors_1
Xsky130_fd_pr__pfet_01v8_4RPJ49_1 gnd vdd vdd gnd gnd vdd vdd vdd gnd vdd gnd gnd
+ vdd gnd gnd gnd vdd vdd vdd vdd gnd vdd gnd gnd gnd gnd gnd gnd gnd vdd gnd vdd
+ gnd gnd vdd gnd gnd vdd vdd gnd vdd gnd gnd vdd gnd gnd vdd vdd gnd gnd vdd vdd
+ vdd gnd gnd vdd vdd gnd gnd vdd vdd gnd vdd gnd vdd gnd gnd gnd vdd gnd gnd gnd
+ vdd vdd gnd gnd vdd vdd gnd gnd vdd vdd gnd gnd gnd vdd vdd vdd vdd vdd vdd vdd
+ vdd vdd gnd gnd vdd vdd vdd gnd vdd vdd vdd vdd vdd gnd vdd vdd gnd vdd vdd gnd
+ gnd gnd gnd gnd vdd vdd vdd gnd vdd vdd gnd vdd gnd vdd vdd vdd gnd gnd vdd vdd
+ gnd vdd vdd vdd vdd gnd vdd gnd gnd gnd vdd vdd vdd gnd gnd gnd gnd vdd gnd gnd
+ gnd vdd gnd gnd gnd gnd vdd gnd gnd vdd vdd sky130_fd_pr__pfet_01v8_4RPJ49
Xcapacitors_1_4 input2 vdd vdd clkb vdd vdd vdd in2 gnd capacitors_1
Xcapacitors_1_5 input2 vdd vdd clkb vdd vdd vdd in3 gnd capacitors_1
Xcapacitors_1_6 input1 vdd vdd clk vdd vdd vdd in4 gnd capacitors_1
Xcapacitors_1_7 input1 vdd vdd clk vdd vdd vdd in5 gnd capacitors_1
Xcapacitors_1_8 input1 vdd vdd clk vdd vdd vdd in6 gnd capacitors_1
Xcapacitors_1_9 input1 vdd vdd clk vdd vdd vdd in7 gnd capacitors_1
Xpmos_cp1_0 m1_12659_300# input2 m1_12464_n576# m1_4341_n519# input1 gnd pmos_cp1
Xsky130_fd_pr__nfet_01v8_NJGC8F_0 vdd gnd gnd vdd vdd gnd gnd vdd gnd vdd gnd gnd
+ vdd gnd gnd gnd vdd gnd vdd vdd gnd vdd vdd vdd vdd gnd vdd vdd gnd vdd vdd gnd
+ gnd gnd gnd gnd vdd gnd gnd vdd gnd gnd gnd vdd gnd gnd vdd gnd gnd gnd vdd vdd
+ gnd gnd vdd gnd gnd vdd gnd gnd gnd vdd vdd vdd gnd gnd gnd gnd vdd gnd vdd gnd
+ vdd gnd gnd vdd gnd vdd vdd vdd vdd vdd vdd gnd gnd gnd gnd gnd vdd gnd gnd vdd
+ vdd gnd vdd vdd vdd vdd gnd vdd gnd gnd gnd gnd gnd vdd vdd vdd vdd gnd vdd vdd
+ vdd vdd gnd vdd gnd vdd vdd gnd gnd vdd gnd gnd vdd vdd vdd gnd gnd vdd gnd gnd
+ gnd vdd vdd gnd vdd vdd vdd gnd vdd vdd gnd gnd gnd vdd vdd vdd gnd vdd vdd vdd
+ vdd vdd vdd gnd vdd gnd vdd gnd gnd gnd sky130_fd_pr__nfet_01v8_NJGC8F
Xcapacitors_1_10 input2 vdd vdd clkb vdd vdd vdd in7 gnd capacitors_1
Xcapacitors_1_11 input2 vdd vdd clkb vdd vdd vdd in6 gnd capacitors_1
Xsky130_fd_pr__nfet_01v8_NJGC8F_1 vdd gnd gnd vdd vdd gnd gnd vdd gnd vdd gnd gnd
+ vdd gnd gnd gnd vdd gnd vdd vdd gnd vdd vdd vdd vdd gnd vdd vdd gnd vdd vdd gnd
+ gnd gnd gnd gnd vdd gnd gnd vdd gnd gnd gnd vdd gnd gnd vdd gnd gnd gnd vdd vdd
+ gnd gnd vdd gnd gnd vdd gnd gnd gnd vdd vdd vdd gnd gnd gnd gnd vdd gnd vdd gnd
+ vdd gnd gnd vdd gnd vdd vdd vdd vdd vdd vdd gnd gnd gnd gnd gnd vdd gnd gnd vdd
+ vdd gnd vdd vdd vdd vdd gnd vdd gnd gnd gnd gnd gnd vdd vdd vdd vdd gnd vdd vdd
+ vdd vdd gnd vdd gnd vdd vdd gnd gnd vdd gnd gnd vdd vdd vdd gnd gnd vdd gnd gnd
+ gnd vdd vdd gnd vdd vdd vdd gnd vdd vdd gnd gnd gnd vdd vdd vdd gnd vdd vdd vdd
+ vdd vdd vdd gnd vdd gnd vdd gnd gnd gnd sky130_fd_pr__nfet_01v8_NJGC8F
Xcapacitors_1_13 input2 vdd vdd clkb vdd vdd vdd in4 gnd capacitors_1
Xcapacitors_1_12 input2 vdd vdd clkb vdd vdd vdd in5 gnd capacitors_1
Xsky130_fd_pr__cap_mim_m3_1_MH6KF8_0 clkb input2 gnd sky130_fd_pr__cap_mim_m3_1_MH6KF8
Xsky130_fd_pr__cap_mim_m3_1_MH6KF8_1 clk input1 gnd sky130_fd_pr__cap_mim_m3_1_MH6KF8
Xsky130_fd_pr__cap_mim_m3_1_MH6KF8_3 m1_12659_300# clkb gnd sky130_fd_pr__cap_mim_m3_1_MH6KF8
Xsky130_fd_pr__cap_mim_m3_1_MH6KF8_2 m1_4341_n519# clk gnd sky130_fd_pr__cap_mim_m3_1_MH6KF8
C0 vin vdd 9.14f
C1 input1 vdd 26.8f
C2 input2 input1 3.06f
C3 vdd clkb 26.2f
C4 m1_12464_n576# clkb 2.21f
C5 clk vdd 32.2f
C6 m1_12464_n576# clk 2.31f
C7 vin clk 2.19f
C8 input2 vdd 26.5f
C9 input1 gnd 31f
C10 input2 gnd 31.1f
C11 capacitors_1_12/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# gnd 2.4f
C12 capacitors_1_12/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# gnd 10.1f
C13 capacitors_1_12/capacitor_8_0/capacitor_7_0/buffer_digital_0/in gnd 2.63f
C14 capacitors_1_13/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# gnd 2.4f
C15 capacitors_1_13/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# gnd 10.1f
C16 capacitors_1_13/capacitor_8_0/capacitor_7_0/buffer_digital_0/in gnd 2.63f
C17 capacitors_1_11/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# gnd 2.39f
C18 capacitors_1_11/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# gnd 10.1f
C19 capacitors_1_11/capacitor_8_0/capacitor_7_0/buffer_digital_0/in gnd 2.63f
C20 capacitors_1_10/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# gnd 2.4f
C21 capacitors_1_10/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# gnd 10.1f
C22 capacitors_1_10/capacitor_8_0/capacitor_7_0/buffer_digital_0/in gnd 2.63f
C23 m1_4341_n519# gnd 4.1f
C24 m1_12659_300# gnd 2.79f
C25 m1_12464_n576# gnd 5.23f
C26 capacitors_1_9/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# gnd 2.4f
C27 capacitors_1_9/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# gnd 10.1f
C28 capacitors_1_9/capacitor_8_0/capacitor_7_0/buffer_digital_0/in gnd 2.63f
C29 capacitors_1_8/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# gnd 2.39f
C30 capacitors_1_8/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# gnd 10.1f
C31 capacitors_1_8/capacitor_8_0/capacitor_7_0/buffer_digital_0/in gnd 2.63f
C32 capacitors_1_7/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# gnd 2.39f
C33 capacitors_1_7/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# gnd 10.1f
C34 capacitors_1_7/capacitor_8_0/capacitor_7_0/buffer_digital_0/in gnd 2.63f
C35 capacitors_1_6/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# gnd 2.39f
C36 capacitors_1_6/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# gnd 10.1f
C37 capacitors_1_6/capacitor_8_0/capacitor_7_0/buffer_digital_0/in gnd 2.63f
C38 capacitors_1_5/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# gnd 2.4f
C39 capacitors_1_5/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# gnd 10.1f
C40 capacitors_1_5/capacitor_8_0/capacitor_7_0/buffer_digital_0/in gnd 2.63f
C41 capacitors_1_4/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# gnd 2.4f
C42 capacitors_1_4/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# gnd 10.1f
C43 capacitors_1_4/capacitor_8_0/capacitor_7_0/buffer_digital_0/in gnd 2.63f
C44 capacitors_1_3/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# gnd 2.4f
C45 capacitors_1_3/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# gnd 10.1f
C46 capacitors_1_3/capacitor_8_0/capacitor_7_0/buffer_digital_0/in gnd 2.63f
C47 capacitors_1_2/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# gnd 2.39f
C48 capacitors_1_2/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# gnd 10.1f
C49 capacitors_1_2/capacitor_8_0/capacitor_7_0/buffer_digital_0/in gnd 2.63f
C50 capacitors_1_1/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# gnd 2.34f
C51 capacitors_1_1/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# gnd 9.98f
C52 capacitors_1_1/capacitor_8_0/capacitor_7_0/buffer_digital_0/in gnd 2.61f
C53 capacitors_1_0/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# gnd 2.34f
C54 capacitors_1_0/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# gnd 9.98f
C55 capacitors_1_0/capacitor_8_0/capacitor_7_0/buffer_digital_0/in gnd 2.61f
C56 capacitor_8_1/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# gnd 2.39f
C57 clkb gnd 91.9f
C58 capacitor_8_1/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# gnd 10.1f
C59 capacitor_8_1/capacitor_7_0/buffer_digital_0/in gnd 2.64f
C60 capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# gnd 2.4f
C61 clk gnd 91.6f
C62 vdd gnd 0.653p
C63 capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# gnd 10.1f
C64 capacitor_8_0/capacitor_7_0/buffer_digital_0/in gnd 2.64f
C65 clock_0/a_2432_n962# gnd 8.68f **FLOATING
C66 clock_0/a_2020_n482# gnd 2.57f **FLOATING
C67 clock_0/a_344_102# gnd 2.81f
C68 clock_0/a_2402_572# gnd 2.17f
C69 clock_0/a_344_n986# gnd 2.38f
C70 clock_0/a_3246_118# gnd 6.83f
C71 g2 gnd 2.34f
C72 vin gnd 10.4f
.ends

.subckt sky130_fd_pr__nfet_01v8_TKGCLY a_n1425_n130# a_1887_n42# a_1503_n42# a_63_n42#
+ a_15_64# a_2127_64# a_n1281_n42# a_111_n130# a_879_n130# a_1263_n130# a_n417_n42#
+ a_2367_n42# a_2223_n130# a_n1761_n42# a_n1905_64# a_n273_n130# a_255_n42# a_n2241_n42#
+ a_735_n42# a_1599_n42# a_1935_64# a_n2429_n42# a_1215_n42# a_n2193_n130# a_n993_n42#
+ a_n1233_n130# a_n753_64# a_n369_64# a_n129_n42# a_2079_n42# a_n1473_n42# a_n609_n42#
+ a_687_n130# a_1071_n130# a_n1953_n42# a_2031_n130# a_n1521_64# a_n1137_64# a_783_64#
+ a_399_64# a_1839_n130# a_n2289_64# a_1791_n42# a_447_n42# a_927_n42# a_n81_n130#
+ a_2319_64# a_n849_n130# a_n321_n42# a_1407_n42# a_1551_64# a_2271_n42# a_1167_64#
+ a_n1185_n42# a_n801_n42# a_n1041_n130# a_n2001_n130# a_n1665_n42# a_n1809_n130#
+ a_495_n130# a_159_n42# a_n2145_n42# a_1647_n130# a_1983_n42# a_639_n42# a_n945_64#
+ a_1119_n42# a_n897_n42# a_n657_n130# a_n513_n42# a_n1377_n42# a_n1713_64# a_n1329_64#
+ a_975_64# a_n1857_n42# a_351_n42# a_n33_n42# a_n1617_n130# a_831_n42# a_1695_n42#
+ a_n2337_n42# a_1311_n42# a_303_n130# a_1743_64# a_1359_64# a_1455_n130# a_n225_n42#
+ a_2175_n42# a_n561_64# a_n1089_n42# a_n177_64# a_n705_n42# a_n465_n130# a_n1569_n42#
+ a_207_64# a_543_n42# a_591_64# a_n2097_64# a_n2385_n130# VSUBS a_n2049_n42# a_1023_n42#
X0 a_63_n42# a_15_64# a_n33_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X1 a_n2241_n42# a_n2289_64# a_n2337_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X2 a_n2337_n42# a_n2385_n130# a_n2429_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X3 a_n2145_n42# a_n2193_n130# a_n2241_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X4 a_n2049_n42# a_n2097_64# a_n2145_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X5 a_2175_n42# a_2127_64# a_2079_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X6 a_2271_n42# a_2223_n130# a_2175_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X7 a_2079_n42# a_2031_n130# a_1983_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X8 a_2367_n42# a_2319_64# a_2271_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X9 a_927_n42# a_879_n130# a_831_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X10 a_1023_n42# a_975_64# a_927_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X11 a_n1953_n42# a_n2001_n130# a_n2049_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X12 a_n1761_n42# a_n1809_n130# a_n1857_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X13 a_n1665_n42# a_n1713_64# a_n1761_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X14 a_n1857_n42# a_n1905_64# a_n1953_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X15 a_n1569_n42# a_n1617_n130# a_n1665_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X16 a_1215_n42# a_1167_64# a_1119_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X17 a_1311_n42# a_1263_n130# a_1215_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X18 a_1503_n42# a_1455_n130# a_1407_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X19 a_1791_n42# a_1743_64# a_1695_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X20 a_1119_n42# a_1071_n130# a_1023_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X21 a_1407_n42# a_1359_64# a_1311_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X22 a_1599_n42# a_1551_64# a_1503_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X23 a_1695_n42# a_1647_n130# a_1599_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X24 a_1887_n42# a_1839_n130# a_1791_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X25 a_1983_n42# a_1935_64# a_1887_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X26 a_n33_n42# a_n81_n130# a_n129_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X27 a_351_n42# a_303_n130# a_255_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X28 a_159_n42# a_111_n130# a_63_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X29 a_255_n42# a_207_64# a_159_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X30 a_447_n42# a_399_64# a_351_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X31 a_543_n42# a_495_n130# a_447_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X32 a_735_n42# a_687_n130# a_639_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X33 a_831_n42# a_783_64# a_735_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X34 a_639_n42# a_591_64# a_543_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X35 a_n1473_n42# a_n1521_64# a_n1569_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X36 a_n1281_n42# a_n1329_64# a_n1377_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X37 a_n1185_n42# a_n1233_n130# a_n1281_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X38 a_n993_n42# a_n1041_n130# a_n1089_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X39 a_n1377_n42# a_n1425_n130# a_n1473_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X40 a_n1089_n42# a_n1137_64# a_n1185_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X41 a_n321_n42# a_n369_64# a_n417_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X42 a_n801_n42# a_n849_n130# a_n897_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X43 a_n705_n42# a_n753_64# a_n801_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X44 a_n609_n42# a_n657_n130# a_n705_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X45 a_n513_n42# a_n561_64# a_n609_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X46 a_n417_n42# a_n465_n130# a_n513_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X47 a_n225_n42# a_n273_n130# a_n321_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X48 a_n129_n42# a_n177_64# a_n225_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X49 a_n897_n42# a_n945_64# a_n993_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
.ends

.subckt nmos_decap_10 a_n2_210# m1_n10_n42# VSUBS
Xsky130_fd_pr__nfet_01v8_NJGC45_0 m1_n10_n42# a_n2_210# m1_n10_n42# a_n2_210# a_n2_210#
+ m1_n10_n42# m1_n10_n42# a_n2_210# a_n2_210# m1_n10_n42# a_n2_210# m1_n10_n42# m1_n10_n42#
+ m1_n10_n42# m1_n10_n42# m1_n10_n42# a_n2_210# m1_n10_n42# a_n2_210# a_n2_210# a_n2_210#
+ VSUBS sky130_fd_pr__nfet_01v8_NJGC45
C0 a_n2_210# VSUBS 2.33f
.ends

.subckt pmos_decap_10 a_12_230# w_6_4# VSUBS
Xsky130_fd_pr__pfet_01v8_4ZKXAA_0 w_6_4# w_6_4# a_12_230# w_6_4# w_6_4# a_12_230#
+ w_6_4# a_12_230# w_6_4# a_12_230# a_12_230# w_6_4# a_12_230# w_6_4# w_6_4# a_12_230#
+ a_12_230# w_6_4# w_6_4# a_12_230# w_6_4# a_12_230# VSUBS sky130_fd_pr__pfet_01v8_4ZKXAA
.ends

.subckt cp1_buffer1 charge_pump1_0/in8 charge_pump1_0/in4 charge_pump1_0/in3 charge_pump1_0/in5
+ charge_pump1_0/in2 charge_pump1_0/vin charge_pump1_0/in6 clk_out clk_in charge_pump1_0/in1
+ charge_pump1_0/m1_12464_n576# charge_pump1_0/in7 gnd vdd
Xsky130_fd_pr__nfet_01v8_HRDN5X_0 vdd gnd vdd vdd vdd vdd gnd gnd gnd vdd gnd vdd
+ gnd gnd gnd gnd vdd vdd gnd gnd gnd vdd vdd vdd vdd vdd gnd gnd gnd gnd vdd gnd
+ sky130_fd_pr__nfet_01v8_HRDN5X
Xcharge_pump1_0 clk_out charge_pump1_0/input1 charge_pump1_0/input2 charge_pump1_0/in1
+ charge_pump1_0/in2 charge_pump1_0/in6 charge_pump1_0/in7 charge_pump1_0/g1 charge_pump1_0/g2
+ charge_pump1_0/clk charge_pump1_0/clkb charge_pump1_0/m1_12464_n576# gnd charge_pump1_0/in4
+ charge_pump1_0/in3 charge_pump1_0/in5 charge_pump1_0/in8 charge_pump1_0/vin vdd
+ gnd charge_pump1
Xsky130_fd_pr__nfet_01v8_TKGCLY_0 vdd gnd gnd gnd vdd vdd gnd vdd vdd vdd gnd gnd
+ vdd gnd vdd vdd gnd gnd gnd gnd vdd gnd gnd vdd gnd vdd vdd vdd gnd gnd gnd gnd
+ vdd vdd gnd vdd vdd vdd vdd vdd vdd vdd gnd gnd gnd vdd vdd vdd gnd gnd vdd gnd
+ vdd gnd gnd vdd vdd gnd vdd vdd gnd gnd vdd gnd gnd vdd gnd gnd vdd gnd gnd vdd
+ vdd vdd gnd gnd gnd vdd gnd gnd gnd gnd vdd vdd vdd vdd gnd gnd vdd gnd vdd gnd
+ vdd gnd vdd gnd vdd vdd vdd gnd gnd gnd sky130_fd_pr__nfet_01v8_TKGCLY
Xbuffer_digital_0 clk_int clk_out vdd gnd buffer_digital
Xbuffer_digital_1 clk_in clk_int vdd gnd buffer_digital
Xnmos_decap_10_0 vdd gnd gnd nmos_decap_10
Xnmos_decap_10_1 vdd gnd gnd nmos_decap_10
Xnmos_decap_10_2 vdd gnd gnd nmos_decap_10
Xnmos_decap_10_3 vdd gnd gnd nmos_decap_10
Xnmos_decap_10_4 vdd gnd gnd nmos_decap_10
Xnmos_decap_10_6 vdd gnd gnd nmos_decap_10
Xnmos_decap_10_5 vdd gnd gnd nmos_decap_10
Xpmos_decap_10_0 gnd vdd gnd pmos_decap_10
Xpmos_decap_10_1 gnd vdd gnd pmos_decap_10
Xpmos_decap_10_2 gnd vdd gnd pmos_decap_10
Xpmos_decap_10_3 gnd vdd gnd pmos_decap_10
Xpmos_decap_10_4 gnd vdd gnd pmos_decap_10
Xpmos_decap_10_5 gnd vdd gnd pmos_decap_10
Xpmos_decap_10_6 gnd vdd gnd pmos_decap_10
Xpmos_decap_10_7 gnd vdd gnd pmos_decap_10
Xpmos_decap_10_9 gnd vdd gnd pmos_decap_10
Xpmos_decap_10_8 gnd vdd gnd pmos_decap_10
C0 vdd clk_out 5.29f
C1 clk_in gnd 6.71f
C2 clk_out gnd 13.1f
C3 charge_pump1_0/input1 gnd 22.5f
C4 charge_pump1_0/input2 gnd 22.2f
C5 charge_pump1_0/capacitors_1_12/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# gnd 2.34f
C6 charge_pump1_0/capacitors_1_12/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# gnd 9.98f
C7 charge_pump1_0/capacitors_1_12/capacitor_8_0/capacitor_7_0/buffer_digital_0/in gnd 2.61f
C8 charge_pump1_0/capacitors_1_13/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# gnd 2.34f
C9 charge_pump1_0/capacitors_1_13/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# gnd 9.98f
C10 charge_pump1_0/capacitors_1_13/capacitor_8_0/capacitor_7_0/buffer_digital_0/in gnd 2.61f
C11 charge_pump1_0/capacitors_1_11/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# gnd 2.34f
C12 charge_pump1_0/capacitors_1_11/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# gnd 9.98f
C13 charge_pump1_0/capacitors_1_11/capacitor_8_0/capacitor_7_0/buffer_digital_0/in gnd 2.61f
C14 charge_pump1_0/capacitors_1_10/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# gnd 2.34f
C15 charge_pump1_0/capacitors_1_10/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# gnd 9.98f
C16 charge_pump1_0/capacitors_1_10/capacitor_8_0/capacitor_7_0/buffer_digital_0/in gnd 2.61f
C17 charge_pump1_0/m1_4341_n519# gnd 3.77f
C18 charge_pump1_0/m1_12659_300# gnd 2.54f
C19 charge_pump1_0/m1_12464_n576# gnd 4.33f
C20 charge_pump1_0/capacitors_1_9/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# gnd 2.34f
C21 charge_pump1_0/capacitors_1_9/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# gnd 9.98f
C22 charge_pump1_0/capacitors_1_9/capacitor_8_0/capacitor_7_0/buffer_digital_0/in gnd 2.61f
C23 charge_pump1_0/capacitors_1_8/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# gnd 2.34f
C24 charge_pump1_0/capacitors_1_8/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# gnd 9.98f
C25 charge_pump1_0/capacitors_1_8/capacitor_8_0/capacitor_7_0/buffer_digital_0/in gnd 2.61f
C26 charge_pump1_0/capacitors_1_7/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# gnd 2.34f
C27 charge_pump1_0/capacitors_1_7/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# gnd 9.98f
C28 charge_pump1_0/capacitors_1_7/capacitor_8_0/capacitor_7_0/buffer_digital_0/in gnd 2.61f
C29 charge_pump1_0/capacitors_1_6/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# gnd 2.34f
C30 charge_pump1_0/capacitors_1_6/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# gnd 9.98f
C31 charge_pump1_0/capacitors_1_6/capacitor_8_0/capacitor_7_0/buffer_digital_0/in gnd 2.61f
C32 charge_pump1_0/capacitors_1_5/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# gnd 2.34f
C33 charge_pump1_0/capacitors_1_5/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# gnd 9.98f
C34 charge_pump1_0/capacitors_1_5/capacitor_8_0/capacitor_7_0/buffer_digital_0/in gnd 2.61f
C35 charge_pump1_0/capacitors_1_4/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# gnd 2.34f
C36 charge_pump1_0/capacitors_1_4/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# gnd 9.98f
C37 charge_pump1_0/capacitors_1_4/capacitor_8_0/capacitor_7_0/buffer_digital_0/in gnd 2.61f
C38 charge_pump1_0/capacitors_1_3/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# gnd 2.34f
C39 charge_pump1_0/capacitors_1_3/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# gnd 9.98f
C40 charge_pump1_0/capacitors_1_3/capacitor_8_0/capacitor_7_0/buffer_digital_0/in gnd 2.61f
C41 charge_pump1_0/capacitors_1_2/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# gnd 2.34f
C42 charge_pump1_0/capacitors_1_2/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# gnd 9.98f
C43 charge_pump1_0/capacitors_1_2/capacitor_8_0/capacitor_7_0/buffer_digital_0/in gnd 2.61f
C44 charge_pump1_0/capacitors_1_1/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# gnd 2.34f
C45 charge_pump1_0/capacitors_1_1/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# gnd 9.98f
C46 charge_pump1_0/capacitors_1_1/capacitor_8_0/capacitor_7_0/buffer_digital_0/in gnd 2.61f
C47 charge_pump1_0/capacitors_1_0/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# gnd 2.34f
C48 charge_pump1_0/capacitors_1_0/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# gnd 9.98f
C49 charge_pump1_0/capacitors_1_0/capacitor_8_0/capacitor_7_0/buffer_digital_0/in gnd 2.61f
C50 charge_pump1_0/capacitor_8_1/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# gnd 2.34f
C51 charge_pump1_0/clkb gnd 90f
C52 charge_pump1_0/capacitor_8_1/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# gnd 9.98f
C53 charge_pump1_0/capacitor_8_1/capacitor_7_0/buffer_digital_0/in gnd 2.61f
C54 charge_pump1_0/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# gnd 2.34f
C55 charge_pump1_0/clk gnd 89.6f
C56 vdd gnd 0.575p
C57 charge_pump1_0/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# gnd 9.98f
C58 charge_pump1_0/capacitor_8_0/capacitor_7_0/buffer_digital_0/in gnd 2.61f
C59 charge_pump1_0/clock_0/a_2432_n962# gnd 8.68f **FLOATING
C60 charge_pump1_0/clock_0/a_2020_n482# gnd 2.57f **FLOATING
C61 charge_pump1_0/clock_0/a_344_102# gnd 2.81f
C62 charge_pump1_0/clock_0/a_2402_572# gnd 2.17f
C63 charge_pump1_0/clock_0/a_344_n986# gnd 2.38f
C64 charge_pump1_0/clock_0/a_3246_118# gnd 6.83f
C65 charge_pump1_0/g2 gnd 2.34f
C66 charge_pump1_0/vin gnd 10.4f
.ends

.subckt charge_pump1_reverse input1 input2 in1 in2 in6 in7 vdd m1_12464_n576# clock_1/clk_in
+ a_3340_18086# in4 in3 in5 gnd in8 nmos_dnw3_0/vs
Xsky130_fd_pr__cap_mim_m3_1_MH6KF8_4 nmos_dnw3_0/clk clock_1/clkb gnd sky130_fd_pr__cap_mim_m3_1_MH6KF8
Xsky130_fd_pr__cap_mim_m3_1_MH6KF8_5 nmos_dnw3_0/clkb clock_1/clk gnd sky130_fd_pr__cap_mim_m3_1_MH6KF8
Xnmos_dnw3_0 nmos_dnw3_0/vs input1 input2 nmos_dnw3_0/clk nmos_dnw3_0/clkb nmos_dnw3_0/vs
+ gnd nmos_dnw3
Xclock_1 clock_1/clk_in vdd gnd clock_1/clk clock_1/clkb clock
Xcapacitor_8_0 vdd input1 clock_1/clkb vdd vdd vdd vdd gnd in8 capacitor_8
Xcapacitor_8_1 vdd input2 clock_1/clk vdd vdd vdd vdd gnd in8 capacitor_8
Xcapacitors_1_0 input1 vdd vdd clock_1/clkb vdd vdd vdd in1 gnd capacitors_1
Xcapacitors_1_1 input2 vdd vdd clock_1/clk vdd vdd vdd in1 gnd capacitors_1
Xcapacitors_1_2 input1 vdd vdd clock_1/clkb vdd vdd vdd in2 gnd capacitors_1
Xsky130_fd_pr__pfet_01v8_4RPJ49_0 gnd vdd vdd gnd gnd vdd vdd vdd gnd vdd gnd gnd
+ vdd gnd gnd gnd vdd vdd vdd vdd gnd vdd gnd gnd gnd gnd gnd gnd gnd vdd gnd vdd
+ gnd gnd vdd gnd gnd vdd vdd gnd vdd gnd gnd vdd gnd gnd vdd vdd gnd gnd vdd vdd
+ vdd gnd gnd vdd vdd gnd gnd vdd vdd gnd vdd gnd vdd gnd gnd gnd vdd gnd gnd gnd
+ vdd vdd gnd gnd vdd vdd gnd gnd vdd vdd gnd gnd gnd vdd vdd vdd vdd vdd vdd vdd
+ vdd vdd gnd gnd vdd vdd vdd gnd vdd vdd vdd vdd vdd gnd vdd vdd gnd vdd vdd gnd
+ gnd gnd gnd gnd vdd vdd vdd gnd vdd vdd gnd vdd gnd vdd vdd vdd gnd gnd vdd vdd
+ gnd vdd vdd vdd vdd gnd vdd gnd gnd gnd vdd vdd vdd gnd gnd gnd gnd vdd gnd gnd
+ gnd vdd gnd gnd gnd gnd vdd gnd gnd vdd vdd sky130_fd_pr__pfet_01v8_4RPJ49
Xsky130_fd_pr__pfet_01v8_4RPJ49_1 gnd vdd vdd gnd gnd vdd vdd vdd gnd vdd gnd gnd
+ vdd gnd gnd gnd vdd vdd vdd vdd gnd vdd gnd gnd gnd gnd gnd gnd gnd vdd gnd vdd
+ gnd gnd vdd gnd gnd vdd vdd gnd vdd gnd gnd vdd gnd gnd vdd vdd gnd gnd vdd vdd
+ vdd gnd gnd vdd vdd gnd gnd vdd vdd gnd vdd gnd vdd gnd gnd gnd vdd gnd gnd gnd
+ vdd vdd gnd gnd vdd vdd gnd gnd vdd vdd gnd gnd gnd vdd vdd vdd vdd vdd vdd vdd
+ vdd vdd gnd gnd vdd vdd vdd gnd vdd vdd vdd vdd vdd gnd vdd vdd gnd vdd vdd gnd
+ gnd gnd gnd gnd vdd vdd vdd gnd vdd vdd gnd vdd gnd vdd vdd vdd gnd gnd vdd vdd
+ gnd vdd vdd vdd vdd gnd vdd gnd gnd gnd vdd vdd vdd gnd gnd gnd gnd vdd gnd gnd
+ gnd vdd gnd gnd gnd gnd vdd gnd gnd vdd vdd sky130_fd_pr__pfet_01v8_4RPJ49
Xcapacitors_1_3 input1 vdd vdd clock_1/clkb vdd vdd vdd in3 gnd capacitors_1
Xcapacitors_1_4 input2 vdd vdd clock_1/clk vdd vdd vdd in2 gnd capacitors_1
Xcapacitors_1_5 input2 vdd vdd clock_1/clk vdd vdd vdd in3 gnd capacitors_1
Xcapacitors_1_6 input1 vdd vdd clock_1/clkb vdd vdd vdd in4 gnd capacitors_1
Xcapacitors_1_7 input1 vdd vdd clock_1/clkb vdd vdd vdd in5 gnd capacitors_1
Xcapacitors_1_8 input1 vdd vdd clock_1/clkb vdd vdd vdd in6 gnd capacitors_1
Xcapacitors_1_9 input1 vdd vdd clock_1/clkb vdd vdd vdd in7 gnd capacitors_1
Xpmos_cp1_0 m1_12659_300# input2 m1_12464_n576# m1_4341_n519# input1 gnd pmos_cp1
Xsky130_fd_pr__nfet_01v8_NJGC8F_0 vdd gnd gnd vdd vdd gnd gnd vdd gnd vdd gnd gnd
+ vdd gnd gnd gnd vdd gnd vdd vdd gnd vdd vdd vdd vdd gnd vdd vdd gnd vdd vdd gnd
+ gnd gnd gnd gnd vdd gnd gnd vdd gnd gnd gnd vdd gnd gnd vdd gnd gnd gnd vdd vdd
+ gnd gnd vdd gnd gnd vdd gnd gnd gnd vdd vdd vdd gnd gnd gnd gnd vdd gnd vdd gnd
+ vdd gnd gnd vdd gnd vdd vdd vdd vdd vdd vdd gnd gnd gnd gnd gnd vdd gnd gnd vdd
+ vdd gnd vdd vdd vdd vdd gnd vdd gnd gnd gnd gnd gnd vdd vdd vdd vdd gnd vdd vdd
+ vdd vdd gnd vdd gnd vdd vdd gnd gnd vdd gnd gnd vdd vdd vdd gnd gnd vdd gnd gnd
+ gnd vdd vdd gnd vdd vdd vdd gnd vdd vdd gnd gnd gnd vdd vdd vdd gnd vdd vdd vdd
+ vdd vdd vdd gnd vdd gnd vdd gnd gnd gnd sky130_fd_pr__nfet_01v8_NJGC8F
Xcapacitors_1_10 input2 vdd vdd clock_1/clk vdd vdd vdd in7 gnd capacitors_1
Xcapacitors_1_11 input2 vdd vdd clock_1/clk vdd vdd vdd in6 gnd capacitors_1
Xsky130_fd_pr__nfet_01v8_NJGC8F_1 vdd gnd gnd vdd vdd gnd gnd vdd gnd vdd gnd gnd
+ vdd gnd gnd gnd vdd gnd vdd vdd gnd vdd vdd vdd vdd gnd vdd vdd gnd vdd vdd gnd
+ gnd gnd gnd gnd vdd gnd gnd vdd gnd gnd gnd vdd gnd gnd vdd gnd gnd gnd vdd vdd
+ gnd gnd vdd gnd gnd vdd gnd gnd gnd vdd vdd vdd gnd gnd gnd gnd vdd gnd vdd gnd
+ vdd gnd gnd vdd gnd vdd vdd vdd vdd vdd vdd gnd gnd gnd gnd gnd vdd gnd gnd vdd
+ vdd gnd vdd vdd vdd vdd gnd vdd gnd gnd gnd gnd gnd vdd vdd vdd vdd gnd vdd vdd
+ vdd vdd gnd vdd gnd vdd vdd gnd gnd vdd gnd gnd vdd vdd vdd gnd gnd vdd gnd gnd
+ gnd vdd vdd gnd vdd vdd vdd gnd vdd vdd gnd gnd gnd vdd vdd vdd gnd vdd vdd vdd
+ vdd vdd vdd gnd vdd gnd vdd gnd gnd gnd sky130_fd_pr__nfet_01v8_NJGC8F
Xcapacitors_1_13 input2 vdd vdd clock_1/clk vdd vdd vdd in4 gnd capacitors_1
Xcapacitors_1_12 input2 vdd vdd clock_1/clk vdd vdd vdd in5 gnd capacitors_1
Xsky130_fd_pr__cap_mim_m3_1_MH6KF8_0 clock_1/clk input2 gnd sky130_fd_pr__cap_mim_m3_1_MH6KF8
Xsky130_fd_pr__cap_mim_m3_1_MH6KF8_1 clock_1/clkb input1 gnd sky130_fd_pr__cap_mim_m3_1_MH6KF8
Xsky130_fd_pr__cap_mim_m3_1_MH6KF8_3 m1_12659_300# clock_1/clk gnd sky130_fd_pr__cap_mim_m3_1_MH6KF8
Xsky130_fd_pr__cap_mim_m3_1_MH6KF8_2 m1_4341_n519# clock_1/clkb gnd sky130_fd_pr__cap_mim_m3_1_MH6KF8
C0 vdd clock_1/clk 28.7f
C1 input2 input1 3.06f
C2 nmos_dnw3_0/vs clock_1/clkb 2.22f
C3 input2 vdd 26.5f
C4 nmos_dnw3_0/vs vdd 9.24f
C5 m1_12464_n576# clock_1/clkb 2.3f
C6 m1_12464_n576# clock_1/clk 2.14f
C7 vdd clock_1/clkb 32.3f
C8 input1 vdd 26.5f
C9 input1 gnd 31.2f
C10 capacitors_1_12/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# gnd 2.4f
C11 capacitors_1_12/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# gnd 10.1f
C12 capacitors_1_12/capacitor_8_0/capacitor_7_0/buffer_digital_0/in gnd 2.63f
C13 capacitors_1_13/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# gnd 2.4f
C14 capacitors_1_13/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# gnd 10.1f
C15 capacitors_1_13/capacitor_8_0/capacitor_7_0/buffer_digital_0/in gnd 2.63f
C16 capacitors_1_11/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# gnd 2.39f
C17 capacitors_1_11/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# gnd 10.1f
C18 capacitors_1_11/capacitor_8_0/capacitor_7_0/buffer_digital_0/in gnd 2.63f
C19 capacitors_1_10/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# gnd 2.4f
C20 capacitors_1_10/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# gnd 10.1f
C21 capacitors_1_10/capacitor_8_0/capacitor_7_0/buffer_digital_0/in gnd 2.63f
C22 m1_4341_n519# gnd 3.77f
C23 input2 gnd 30.6f
C24 m1_12659_300# gnd 3.03f
C25 m1_12464_n576# gnd 5.5f
C26 capacitors_1_9/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# gnd 2.4f
C27 capacitors_1_9/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# gnd 10.1f
C28 capacitors_1_9/capacitor_8_0/capacitor_7_0/buffer_digital_0/in gnd 2.63f
C29 capacitors_1_8/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# gnd 2.39f
C30 capacitors_1_8/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# gnd 10.1f
C31 capacitors_1_8/capacitor_8_0/capacitor_7_0/buffer_digital_0/in gnd 2.63f
C32 capacitors_1_7/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# gnd 2.39f
C33 capacitors_1_7/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# gnd 10.1f
C34 capacitors_1_7/capacitor_8_0/capacitor_7_0/buffer_digital_0/in gnd 2.63f
C35 capacitors_1_6/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# gnd 2.39f
C36 capacitors_1_6/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# gnd 10.1f
C37 capacitors_1_6/capacitor_8_0/capacitor_7_0/buffer_digital_0/in gnd 2.63f
C38 capacitors_1_5/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# gnd 2.4f
C39 capacitors_1_5/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# gnd 10.1f
C40 capacitors_1_5/capacitor_8_0/capacitor_7_0/buffer_digital_0/in gnd 2.63f
C41 capacitors_1_4/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# gnd 2.4f
C42 capacitors_1_4/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# gnd 10.1f
C43 capacitors_1_4/capacitor_8_0/capacitor_7_0/buffer_digital_0/in gnd 2.63f
C44 capacitors_1_3/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# gnd 2.4f
C45 capacitors_1_3/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# gnd 10.1f
C46 capacitors_1_3/capacitor_8_0/capacitor_7_0/buffer_digital_0/in gnd 2.63f
C47 capacitors_1_2/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# gnd 2.39f
C48 capacitors_1_2/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# gnd 10.1f
C49 capacitors_1_2/capacitor_8_0/capacitor_7_0/buffer_digital_0/in gnd 2.63f
C50 capacitors_1_1/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# gnd 2.34f
C51 capacitors_1_1/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# gnd 9.98f
C52 capacitors_1_1/capacitor_8_0/capacitor_7_0/buffer_digital_0/in gnd 2.61f
C53 capacitors_1_0/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# gnd 2.34f
C54 capacitors_1_0/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# gnd 9.98f
C55 capacitors_1_0/capacitor_8_0/capacitor_7_0/buffer_digital_0/in gnd 2.61f
C56 capacitor_8_1/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# gnd 2.39f
C57 clock_1/clk gnd 96.8f
C58 capacitor_8_1/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# gnd 10.1f
C59 capacitor_8_1/capacitor_7_0/buffer_digital_0/in gnd 2.64f
C60 capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# gnd 2.4f
C61 clock_1/clkb gnd 0.105p
C62 vdd gnd 0.66p
C63 capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# gnd 10.1f
C64 capacitor_8_0/capacitor_7_0/buffer_digital_0/in gnd 2.64f
C65 clock_1/a_2432_n962# gnd 8.69f **FLOATING
C66 clock_1/a_2020_n482# gnd 2.57f **FLOATING
C67 clock_1/a_344_102# gnd 2.81f
C68 clock_1/a_2402_572# gnd 2.17f
C69 clock_1/a_344_n986# gnd 2.38f
C70 clock_1/a_3246_118# gnd 6.83f
C71 nmos_dnw3_0/vs gnd 10.4f
.ends

.subckt cp1_buffer1_reverse charge_pump1_reverse_0/m1_12464_n576# charge_pump1_reverse_0/in6
+ charge_pump1_reverse_0/in7 charge_pump1_reverse_0/in1 buffer_digital_0/in charge_pump1_reverse_0/in8
+ buffer_digital_1/VDD charge_pump1_reverse_0/nmos_dnw3_0/vs charge_pump1_reverse_0/in4
+ charge_pump1_reverse_0/in3 buffer_digital_1/i charge_pump1_reverse_0/in5 charge_pump1_reverse_0/in2
+ VSUBS
Xpmos_decap_10_10 VSUBS buffer_digital_1/VDD VSUBS pmos_decap_10
Xpmos_decap_10_11 VSUBS buffer_digital_1/VDD VSUBS pmos_decap_10
Xpmos_decap_10_12 VSUBS buffer_digital_1/VDD VSUBS pmos_decap_10
Xpmos_decap_10_13 VSUBS buffer_digital_1/VDD VSUBS pmos_decap_10
Xpmos_decap_10_14 VSUBS buffer_digital_1/VDD VSUBS pmos_decap_10
Xcharge_pump1_reverse_0 charge_pump1_reverse_0/input1 charge_pump1_reverse_0/input2
+ charge_pump1_reverse_0/in1 charge_pump1_reverse_0/in2 charge_pump1_reverse_0/in6
+ charge_pump1_reverse_0/in7 buffer_digital_1/VDD charge_pump1_reverse_0/m1_12464_n576#
+ buffer_digital_0/in VSUBS charge_pump1_reverse_0/in4 charge_pump1_reverse_0/in3
+ charge_pump1_reverse_0/in5 VSUBS charge_pump1_reverse_0/in8 charge_pump1_reverse_0/nmos_dnw3_0/vs
+ charge_pump1_reverse
Xbuffer_digital_0 buffer_digital_0/i buffer_digital_0/in buffer_digital_1/VDD VSUBS
+ buffer_digital
Xbuffer_digital_1 buffer_digital_1/i buffer_digital_0/i buffer_digital_1/VDD VSUBS
+ buffer_digital
Xnmos_decap_10_0 buffer_digital_1/VDD VSUBS VSUBS nmos_decap_10
Xnmos_decap_10_1 buffer_digital_1/VDD VSUBS VSUBS nmos_decap_10
Xnmos_decap_10_2 buffer_digital_1/VDD VSUBS VSUBS nmos_decap_10
Xnmos_decap_10_3 buffer_digital_1/VDD VSUBS VSUBS nmos_decap_10
Xnmos_decap_10_4 buffer_digital_1/VDD VSUBS VSUBS nmos_decap_10
Xnmos_decap_10_10 buffer_digital_1/VDD VSUBS VSUBS nmos_decap_10
Xnmos_decap_10_11 buffer_digital_1/VDD VSUBS VSUBS nmos_decap_10
Xnmos_decap_10_5 buffer_digital_1/VDD VSUBS VSUBS nmos_decap_10
Xnmos_decap_10_6 buffer_digital_1/VDD VSUBS VSUBS nmos_decap_10
Xnmos_decap_10_12 buffer_digital_1/VDD VSUBS VSUBS nmos_decap_10
Xnmos_decap_10_7 buffer_digital_1/VDD VSUBS VSUBS nmos_decap_10
Xnmos_decap_10_8 buffer_digital_1/VDD VSUBS VSUBS nmos_decap_10
Xpmos_decap_10_0 VSUBS buffer_digital_1/VDD VSUBS pmos_decap_10
Xnmos_decap_10_9 buffer_digital_1/VDD VSUBS VSUBS nmos_decap_10
Xpmos_decap_10_1 VSUBS buffer_digital_1/VDD VSUBS pmos_decap_10
Xpmos_decap_10_2 VSUBS buffer_digital_1/VDD VSUBS pmos_decap_10
Xpmos_decap_10_3 VSUBS buffer_digital_1/VDD VSUBS pmos_decap_10
Xpmos_decap_10_4 VSUBS buffer_digital_1/VDD VSUBS pmos_decap_10
Xpmos_decap_10_5 VSUBS buffer_digital_1/VDD VSUBS pmos_decap_10
Xpmos_decap_10_6 VSUBS buffer_digital_1/VDD VSUBS pmos_decap_10
Xpmos_decap_10_7 VSUBS buffer_digital_1/VDD VSUBS pmos_decap_10
Xpmos_decap_10_9 VSUBS buffer_digital_1/VDD VSUBS pmos_decap_10
Xpmos_decap_10_8 VSUBS buffer_digital_1/VDD VSUBS pmos_decap_10
C0 charge_pump1_reverse_0/clock_1/clkb buffer_digital_1/VDD 2.74f
C1 buffer_digital_0/in buffer_digital_1/VDD 5.98f
C2 buffer_digital_1/i VSUBS 6.66f
C3 charge_pump1_reverse_0/input1 VSUBS 22.6f
C4 charge_pump1_reverse_0/capacitors_1_12/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# VSUBS 2.34f
C5 charge_pump1_reverse_0/capacitors_1_12/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# VSUBS 9.98f
C6 charge_pump1_reverse_0/capacitors_1_12/capacitor_8_0/capacitor_7_0/buffer_digital_0/in VSUBS 2.61f
C7 charge_pump1_reverse_0/capacitors_1_13/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# VSUBS 2.34f
C8 charge_pump1_reverse_0/capacitors_1_13/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# VSUBS 9.98f
C9 charge_pump1_reverse_0/capacitors_1_13/capacitor_8_0/capacitor_7_0/buffer_digital_0/in VSUBS 2.61f
C10 charge_pump1_reverse_0/capacitors_1_11/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# VSUBS 2.34f
C11 charge_pump1_reverse_0/capacitors_1_11/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# VSUBS 9.98f
C12 charge_pump1_reverse_0/capacitors_1_11/capacitor_8_0/capacitor_7_0/buffer_digital_0/in VSUBS 2.61f
C13 charge_pump1_reverse_0/capacitors_1_10/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# VSUBS 2.34f
C14 charge_pump1_reverse_0/capacitors_1_10/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# VSUBS 9.98f
C15 charge_pump1_reverse_0/capacitors_1_10/capacitor_8_0/capacitor_7_0/buffer_digital_0/in VSUBS 2.61f
C16 charge_pump1_reverse_0/m1_4341_n519# VSUBS 3.33f
C17 charge_pump1_reverse_0/input2 VSUBS 22.2f
C18 charge_pump1_reverse_0/m1_12659_300# VSUBS 2.68f
C19 charge_pump1_reverse_0/m1_12464_n576# VSUBS 4.64f
C20 charge_pump1_reverse_0/capacitors_1_9/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# VSUBS 2.34f
C21 charge_pump1_reverse_0/capacitors_1_9/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# VSUBS 9.98f
C22 charge_pump1_reverse_0/capacitors_1_9/capacitor_8_0/capacitor_7_0/buffer_digital_0/in VSUBS 2.61f
C23 charge_pump1_reverse_0/capacitors_1_8/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# VSUBS 2.34f
C24 charge_pump1_reverse_0/capacitors_1_8/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# VSUBS 9.98f
C25 charge_pump1_reverse_0/capacitors_1_8/capacitor_8_0/capacitor_7_0/buffer_digital_0/in VSUBS 2.61f
C26 charge_pump1_reverse_0/capacitors_1_7/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# VSUBS 2.34f
C27 charge_pump1_reverse_0/capacitors_1_7/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# VSUBS 9.98f
C28 charge_pump1_reverse_0/capacitors_1_7/capacitor_8_0/capacitor_7_0/buffer_digital_0/in VSUBS 2.61f
C29 charge_pump1_reverse_0/capacitors_1_6/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# VSUBS 2.34f
C30 charge_pump1_reverse_0/capacitors_1_6/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# VSUBS 9.98f
C31 charge_pump1_reverse_0/capacitors_1_6/capacitor_8_0/capacitor_7_0/buffer_digital_0/in VSUBS 2.61f
C32 charge_pump1_reverse_0/capacitors_1_5/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# VSUBS 2.34f
C33 charge_pump1_reverse_0/capacitors_1_5/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# VSUBS 9.98f
C34 charge_pump1_reverse_0/capacitors_1_5/capacitor_8_0/capacitor_7_0/buffer_digital_0/in VSUBS 2.61f
C35 charge_pump1_reverse_0/capacitors_1_4/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# VSUBS 2.34f
C36 charge_pump1_reverse_0/capacitors_1_4/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# VSUBS 9.98f
C37 charge_pump1_reverse_0/capacitors_1_4/capacitor_8_0/capacitor_7_0/buffer_digital_0/in VSUBS 2.61f
C38 charge_pump1_reverse_0/capacitors_1_3/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# VSUBS 2.34f
C39 charge_pump1_reverse_0/capacitors_1_3/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# VSUBS 9.98f
C40 charge_pump1_reverse_0/capacitors_1_3/capacitor_8_0/capacitor_7_0/buffer_digital_0/in VSUBS 2.61f
C41 charge_pump1_reverse_0/capacitors_1_2/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# VSUBS 2.34f
C42 charge_pump1_reverse_0/capacitors_1_2/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# VSUBS 9.98f
C43 charge_pump1_reverse_0/capacitors_1_2/capacitor_8_0/capacitor_7_0/buffer_digital_0/in VSUBS 2.61f
C44 charge_pump1_reverse_0/capacitors_1_1/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# VSUBS 2.34f
C45 charge_pump1_reverse_0/capacitors_1_1/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# VSUBS 9.98f
C46 charge_pump1_reverse_0/capacitors_1_1/capacitor_8_0/capacitor_7_0/buffer_digital_0/in VSUBS 2.61f
C47 charge_pump1_reverse_0/capacitors_1_0/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# VSUBS 2.34f
C48 charge_pump1_reverse_0/capacitors_1_0/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# VSUBS 9.98f
C49 charge_pump1_reverse_0/capacitors_1_0/capacitor_8_0/capacitor_7_0/buffer_digital_0/in VSUBS 2.61f
C50 charge_pump1_reverse_0/capacitor_8_1/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# VSUBS 2.34f
C51 charge_pump1_reverse_0/clock_1/clk VSUBS 94.7f
C52 charge_pump1_reverse_0/capacitor_8_1/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# VSUBS 9.98f
C53 charge_pump1_reverse_0/capacitor_8_1/capacitor_7_0/buffer_digital_0/in VSUBS 2.61f
C54 charge_pump1_reverse_0/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# VSUBS 2.34f
C55 charge_pump1_reverse_0/clock_1/clkb VSUBS 0.101p
C56 buffer_digital_1/VDD VSUBS 0.575p
C57 charge_pump1_reverse_0/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# VSUBS 9.98f
C58 charge_pump1_reverse_0/capacitor_8_0/capacitor_7_0/buffer_digital_0/in VSUBS 2.61f
C59 charge_pump1_reverse_0/clock_1/a_2432_n962# VSUBS 8.68f **FLOATING
C60 charge_pump1_reverse_0/clock_1/a_2020_n482# VSUBS 2.57f **FLOATING
C61 charge_pump1_reverse_0/clock_1/a_344_102# VSUBS 2.81f
C62 charge_pump1_reverse_0/clock_1/a_2402_572# VSUBS 2.17f
C63 charge_pump1_reverse_0/clock_1/a_344_n986# VSUBS 2.38f
C64 buffer_digital_0/in VSUBS 16.5f
C65 charge_pump1_reverse_0/clock_1/a_3246_118# VSUBS 6.83f
C66 charge_pump1_reverse_0/nmos_dnw3_0/vs VSUBS 10.3f
.ends

.subckt cp1_buffer_5stage cp1_buffer1_2/charge_pump1_0/in2 cp1_buffer1_2/charge_pump1_0/in8
+ cp1_buffer1_2/charge_pump1_0/in7 cp1_buffer1_2/charge_pump1_0/in6 cp1_buffer1_2/charge_pump1_0/in1
+ cp1_buffer1_2/charge_pump1_0/in5 cp1_buffer1_2/charge_pump1_0/m1_12464_n576# cp1_buffer1_reverse_1/charge_pump1_reverse_0/nmos_dnw3_0/vs
+ cp1_buffer1_0/clk_in cp1_buffer1_2/charge_pump1_0/in4 cp1_buffer1_reverse_0/charge_pump1_reverse_0/nmos_dnw3_0/vs
+ cp1_buffer1_0/charge_pump1_0/vin cp1_buffer1_1/charge_pump1_0/vin cp1_buffer1_2/vdd
+ VSUBS cp1_buffer1_2/charge_pump1_0/in3 cp1_buffer1_2/charge_pump1_0/vin
Xcp1_buffer1_0 cp1_buffer1_2/charge_pump1_0/in8 cp1_buffer1_2/charge_pump1_0/in4 cp1_buffer1_2/charge_pump1_0/in3
+ cp1_buffer1_2/charge_pump1_0/in5 cp1_buffer1_2/charge_pump1_0/in2 cp1_buffer1_0/charge_pump1_0/vin
+ cp1_buffer1_2/charge_pump1_0/in6 cp1_buffer1_0/clk_out cp1_buffer1_0/clk_in cp1_buffer1_2/charge_pump1_0/in1
+ cp1_buffer1_reverse_0/charge_pump1_reverse_0/nmos_dnw3_0/vs cp1_buffer1_2/charge_pump1_0/in7
+ VSUBS cp1_buffer1_2/vdd cp1_buffer1
Xcp1_buffer1_1 cp1_buffer1_2/charge_pump1_0/in8 cp1_buffer1_2/charge_pump1_0/in4 cp1_buffer1_2/charge_pump1_0/in3
+ cp1_buffer1_2/charge_pump1_0/in5 cp1_buffer1_2/charge_pump1_0/in2 cp1_buffer1_1/charge_pump1_0/vin
+ cp1_buffer1_2/charge_pump1_0/in6 cp1_buffer1_1/clk_out cp1_buffer1_1/clk_in cp1_buffer1_2/charge_pump1_0/in1
+ cp1_buffer1_reverse_1/charge_pump1_reverse_0/nmos_dnw3_0/vs cp1_buffer1_2/charge_pump1_0/in7
+ VSUBS cp1_buffer1_2/vdd cp1_buffer1
Xcp1_buffer1_2 cp1_buffer1_2/charge_pump1_0/in8 cp1_buffer1_2/charge_pump1_0/in4 cp1_buffer1_2/charge_pump1_0/in3
+ cp1_buffer1_2/charge_pump1_0/in5 cp1_buffer1_2/charge_pump1_0/in2 cp1_buffer1_2/charge_pump1_0/vin
+ cp1_buffer1_2/charge_pump1_0/in6 cp1_buffer1_2/clk_out cp1_buffer1_2/clk_in cp1_buffer1_2/charge_pump1_0/in1
+ cp1_buffer1_2/charge_pump1_0/m1_12464_n576# cp1_buffer1_2/charge_pump1_0/in7 VSUBS
+ cp1_buffer1_2/vdd cp1_buffer1
Xcp1_buffer1_reverse_0 cp1_buffer1_1/charge_pump1_0/vin cp1_buffer1_2/charge_pump1_0/in3
+ cp1_buffer1_2/charge_pump1_0/in2 cp1_buffer1_2/charge_pump1_0/in8 cp1_buffer1_1/clk_in
+ cp1_buffer1_2/charge_pump1_0/in1 cp1_buffer1_2/vdd cp1_buffer1_reverse_0/charge_pump1_reverse_0/nmos_dnw3_0/vs
+ cp1_buffer1_2/charge_pump1_0/in5 cp1_buffer1_2/charge_pump1_0/in6 cp1_buffer1_0/clk_out
+ cp1_buffer1_2/charge_pump1_0/in4 cp1_buffer1_2/charge_pump1_0/in7 VSUBS cp1_buffer1_reverse
Xcp1_buffer1_reverse_1 cp1_buffer1_2/charge_pump1_0/vin cp1_buffer1_2/charge_pump1_0/in3
+ cp1_buffer1_2/charge_pump1_0/in2 cp1_buffer1_2/charge_pump1_0/in8 cp1_buffer1_2/clk_in
+ cp1_buffer1_2/charge_pump1_0/in1 cp1_buffer1_2/vdd cp1_buffer1_reverse_1/charge_pump1_reverse_0/nmos_dnw3_0/vs
+ cp1_buffer1_2/charge_pump1_0/in5 cp1_buffer1_2/charge_pump1_0/in6 cp1_buffer1_1/clk_out
+ cp1_buffer1_2/charge_pump1_0/in4 cp1_buffer1_2/charge_pump1_0/in7 VSUBS cp1_buffer1_reverse
C0 cp1_buffer1_2/vdd cp1_buffer1_0/clk_out 2.01f
C1 cp1_buffer1_2/vdd cp1_buffer1_2/charge_pump1_0/in4 3.95f
C2 cp1_buffer1_2/vdd cp1_buffer1_2/charge_pump1_0/in3 3.9f
C3 cp1_buffer1_2/vdd cp1_buffer1_2/charge_pump1_0/in1 4f
C4 cp1_buffer1_2/vdd cp1_buffer1_2/charge_pump1_0/in6 4.05f
C5 cp1_buffer1_2/vdd cp1_buffer1_1/clk_out 2.55f
C6 cp1_buffer1_2/vdd cp1_buffer1_2/charge_pump1_0/in2 3.97f
C7 cp1_buffer1_2/vdd cp1_buffer1_2/charge_pump1_0/in7 3.64f
C8 cp1_buffer1_2/vdd cp1_buffer1_2/charge_pump1_0/in5 3.91f
C9 cp1_buffer1_2/vdd cp1_buffer1_2/charge_pump1_0/in8 3.7f
C10 cp1_buffer1_2/vdd cp1_buffer1_1/clk_in 4.13f
C11 cp1_buffer1_reverse_1/charge_pump1_reverse_0/input1 VSUBS 22.6f
C12 cp1_buffer1_reverse_1/charge_pump1_reverse_0/capacitors_1_12/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# VSUBS 2.34f
C13 cp1_buffer1_reverse_1/charge_pump1_reverse_0/capacitors_1_12/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# VSUBS 9.98f
C14 cp1_buffer1_reverse_1/charge_pump1_reverse_0/capacitors_1_12/capacitor_8_0/capacitor_7_0/buffer_digital_0/in VSUBS 2.61f
C15 cp1_buffer1_reverse_1/charge_pump1_reverse_0/capacitors_1_13/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# VSUBS 2.34f
C16 cp1_buffer1_reverse_1/charge_pump1_reverse_0/capacitors_1_13/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# VSUBS 9.98f
C17 cp1_buffer1_reverse_1/charge_pump1_reverse_0/capacitors_1_13/capacitor_8_0/capacitor_7_0/buffer_digital_0/in VSUBS 2.61f
C18 cp1_buffer1_reverse_1/charge_pump1_reverse_0/capacitors_1_11/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# VSUBS 2.34f
C19 cp1_buffer1_reverse_1/charge_pump1_reverse_0/capacitors_1_11/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# VSUBS 9.98f
C20 cp1_buffer1_reverse_1/charge_pump1_reverse_0/capacitors_1_11/capacitor_8_0/capacitor_7_0/buffer_digital_0/in VSUBS 2.61f
C21 cp1_buffer1_reverse_1/charge_pump1_reverse_0/capacitors_1_10/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# VSUBS 2.34f
C22 cp1_buffer1_reverse_1/charge_pump1_reverse_0/capacitors_1_10/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# VSUBS 9.98f
C23 cp1_buffer1_reverse_1/charge_pump1_reverse_0/capacitors_1_10/capacitor_8_0/capacitor_7_0/buffer_digital_0/in VSUBS 2.61f
C24 cp1_buffer1_reverse_1/charge_pump1_reverse_0/m1_4341_n519# VSUBS 3.33f
C25 cp1_buffer1_reverse_1/charge_pump1_reverse_0/input2 VSUBS 22.2f
C26 cp1_buffer1_reverse_1/charge_pump1_reverse_0/m1_12659_300# VSUBS 2.68f
C27 cp1_buffer1_reverse_1/charge_pump1_reverse_0/capacitors_1_9/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# VSUBS 2.34f
C28 cp1_buffer1_reverse_1/charge_pump1_reverse_0/capacitors_1_9/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# VSUBS 9.98f
C29 cp1_buffer1_reverse_1/charge_pump1_reverse_0/capacitors_1_9/capacitor_8_0/capacitor_7_0/buffer_digital_0/in VSUBS 2.61f
C30 cp1_buffer1_reverse_1/charge_pump1_reverse_0/capacitors_1_8/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# VSUBS 2.34f
C31 cp1_buffer1_reverse_1/charge_pump1_reverse_0/capacitors_1_8/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# VSUBS 9.98f
C32 cp1_buffer1_reverse_1/charge_pump1_reverse_0/capacitors_1_8/capacitor_8_0/capacitor_7_0/buffer_digital_0/in VSUBS 2.61f
C33 cp1_buffer1_reverse_1/charge_pump1_reverse_0/capacitors_1_7/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# VSUBS 2.34f
C34 cp1_buffer1_reverse_1/charge_pump1_reverse_0/capacitors_1_7/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# VSUBS 9.98f
C35 cp1_buffer1_reverse_1/charge_pump1_reverse_0/capacitors_1_7/capacitor_8_0/capacitor_7_0/buffer_digital_0/in VSUBS 2.61f
C36 cp1_buffer1_reverse_1/charge_pump1_reverse_0/capacitors_1_6/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# VSUBS 2.34f
C37 cp1_buffer1_reverse_1/charge_pump1_reverse_0/capacitors_1_6/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# VSUBS 9.98f
C38 cp1_buffer1_reverse_1/charge_pump1_reverse_0/capacitors_1_6/capacitor_8_0/capacitor_7_0/buffer_digital_0/in VSUBS 2.61f
C39 cp1_buffer1_reverse_1/charge_pump1_reverse_0/capacitors_1_5/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# VSUBS 2.34f
C40 cp1_buffer1_reverse_1/charge_pump1_reverse_0/capacitors_1_5/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# VSUBS 9.98f
C41 cp1_buffer1_reverse_1/charge_pump1_reverse_0/capacitors_1_5/capacitor_8_0/capacitor_7_0/buffer_digital_0/in VSUBS 2.61f
C42 cp1_buffer1_reverse_1/charge_pump1_reverse_0/capacitors_1_4/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# VSUBS 2.34f
C43 cp1_buffer1_reverse_1/charge_pump1_reverse_0/capacitors_1_4/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# VSUBS 9.98f
C44 cp1_buffer1_reverse_1/charge_pump1_reverse_0/capacitors_1_4/capacitor_8_0/capacitor_7_0/buffer_digital_0/in VSUBS 2.61f
C45 cp1_buffer1_reverse_1/charge_pump1_reverse_0/capacitors_1_3/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# VSUBS 2.34f
C46 cp1_buffer1_reverse_1/charge_pump1_reverse_0/capacitors_1_3/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# VSUBS 9.98f
C47 cp1_buffer1_reverse_1/charge_pump1_reverse_0/capacitors_1_3/capacitor_8_0/capacitor_7_0/buffer_digital_0/in VSUBS 2.61f
C48 cp1_buffer1_reverse_1/charge_pump1_reverse_0/capacitors_1_2/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# VSUBS 2.34f
C49 cp1_buffer1_reverse_1/charge_pump1_reverse_0/capacitors_1_2/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# VSUBS 9.98f
C50 cp1_buffer1_reverse_1/charge_pump1_reverse_0/capacitors_1_2/capacitor_8_0/capacitor_7_0/buffer_digital_0/in VSUBS 2.61f
C51 cp1_buffer1_reverse_1/charge_pump1_reverse_0/capacitors_1_1/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# VSUBS 2.34f
C52 cp1_buffer1_reverse_1/charge_pump1_reverse_0/capacitors_1_1/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# VSUBS 9.98f
C53 cp1_buffer1_reverse_1/charge_pump1_reverse_0/capacitors_1_1/capacitor_8_0/capacitor_7_0/buffer_digital_0/in VSUBS 2.61f
C54 cp1_buffer1_reverse_1/charge_pump1_reverse_0/capacitors_1_0/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# VSUBS 2.34f
C55 cp1_buffer1_reverse_1/charge_pump1_reverse_0/capacitors_1_0/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# VSUBS 9.98f
C56 cp1_buffer1_reverse_1/charge_pump1_reverse_0/capacitors_1_0/capacitor_8_0/capacitor_7_0/buffer_digital_0/in VSUBS 2.61f
C57 cp1_buffer1_2/charge_pump1_0/in8 VSUBS 11.3f
C58 cp1_buffer1_reverse_1/charge_pump1_reverse_0/capacitor_8_1/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# VSUBS 2.34f
C59 cp1_buffer1_reverse_1/charge_pump1_reverse_0/clock_1/clk VSUBS 94.6f
C60 cp1_buffer1_reverse_1/charge_pump1_reverse_0/capacitor_8_1/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# VSUBS 9.98f
C61 cp1_buffer1_reverse_1/charge_pump1_reverse_0/capacitor_8_1/capacitor_7_0/buffer_digital_0/in VSUBS 2.61f
C62 cp1_buffer1_reverse_1/charge_pump1_reverse_0/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# VSUBS 2.34f
C63 cp1_buffer1_reverse_1/charge_pump1_reverse_0/clock_1/clkb VSUBS 0.101p
C64 cp1_buffer1_reverse_1/charge_pump1_reverse_0/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# VSUBS 9.98f
C65 cp1_buffer1_reverse_1/charge_pump1_reverse_0/capacitor_8_0/capacitor_7_0/buffer_digital_0/in VSUBS 2.61f
C66 cp1_buffer1_reverse_1/charge_pump1_reverse_0/clock_1/a_2432_n962# VSUBS 8.68f **FLOATING
C67 cp1_buffer1_reverse_1/charge_pump1_reverse_0/clock_1/a_2020_n482# VSUBS 2.57f **FLOATING
C68 cp1_buffer1_reverse_1/charge_pump1_reverse_0/clock_1/a_344_102# VSUBS 2.81f
C69 cp1_buffer1_reverse_1/charge_pump1_reverse_0/clock_1/a_2402_572# VSUBS 2.17f
C70 cp1_buffer1_reverse_1/charge_pump1_reverse_0/clock_1/a_344_n986# VSUBS 2.38f
C71 cp1_buffer1_2/clk_in VSUBS 7.49f
C72 cp1_buffer1_reverse_1/charge_pump1_reverse_0/clock_1/a_3246_118# VSUBS 6.83f
C73 cp1_buffer1_reverse_0/charge_pump1_reverse_0/input1 VSUBS 22.6f
C74 cp1_buffer1_reverse_0/charge_pump1_reverse_0/capacitors_1_12/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# VSUBS 2.34f
C75 cp1_buffer1_reverse_0/charge_pump1_reverse_0/capacitors_1_12/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# VSUBS 9.98f
C76 cp1_buffer1_reverse_0/charge_pump1_reverse_0/capacitors_1_12/capacitor_8_0/capacitor_7_0/buffer_digital_0/in VSUBS 2.61f
C77 cp1_buffer1_reverse_0/charge_pump1_reverse_0/capacitors_1_13/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# VSUBS 2.34f
C78 cp1_buffer1_reverse_0/charge_pump1_reverse_0/capacitors_1_13/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# VSUBS 9.98f
C79 cp1_buffer1_reverse_0/charge_pump1_reverse_0/capacitors_1_13/capacitor_8_0/capacitor_7_0/buffer_digital_0/in VSUBS 2.61f
C80 cp1_buffer1_reverse_0/charge_pump1_reverse_0/capacitors_1_11/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# VSUBS 2.34f
C81 cp1_buffer1_reverse_0/charge_pump1_reverse_0/capacitors_1_11/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# VSUBS 9.98f
C82 cp1_buffer1_reverse_0/charge_pump1_reverse_0/capacitors_1_11/capacitor_8_0/capacitor_7_0/buffer_digital_0/in VSUBS 2.61f
C83 cp1_buffer1_reverse_0/charge_pump1_reverse_0/capacitors_1_10/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# VSUBS 2.34f
C84 cp1_buffer1_reverse_0/charge_pump1_reverse_0/capacitors_1_10/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# VSUBS 9.98f
C85 cp1_buffer1_reverse_0/charge_pump1_reverse_0/capacitors_1_10/capacitor_8_0/capacitor_7_0/buffer_digital_0/in VSUBS 2.61f
C86 cp1_buffer1_reverse_0/charge_pump1_reverse_0/m1_4341_n519# VSUBS 3.33f
C87 cp1_buffer1_reverse_0/charge_pump1_reverse_0/input2 VSUBS 22.2f
C88 cp1_buffer1_reverse_0/charge_pump1_reverse_0/m1_12659_300# VSUBS 2.68f
C89 cp1_buffer1_reverse_0/charge_pump1_reverse_0/capacitors_1_9/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# VSUBS 2.34f
C90 cp1_buffer1_reverse_0/charge_pump1_reverse_0/capacitors_1_9/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# VSUBS 9.98f
C91 cp1_buffer1_reverse_0/charge_pump1_reverse_0/capacitors_1_9/capacitor_8_0/capacitor_7_0/buffer_digital_0/in VSUBS 2.61f
C92 cp1_buffer1_reverse_0/charge_pump1_reverse_0/capacitors_1_8/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# VSUBS 2.34f
C93 cp1_buffer1_reverse_0/charge_pump1_reverse_0/capacitors_1_8/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# VSUBS 9.98f
C94 cp1_buffer1_reverse_0/charge_pump1_reverse_0/capacitors_1_8/capacitor_8_0/capacitor_7_0/buffer_digital_0/in VSUBS 2.61f
C95 cp1_buffer1_reverse_0/charge_pump1_reverse_0/capacitors_1_7/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# VSUBS 2.34f
C96 cp1_buffer1_reverse_0/charge_pump1_reverse_0/capacitors_1_7/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# VSUBS 9.98f
C97 cp1_buffer1_reverse_0/charge_pump1_reverse_0/capacitors_1_7/capacitor_8_0/capacitor_7_0/buffer_digital_0/in VSUBS 2.61f
C98 cp1_buffer1_reverse_0/charge_pump1_reverse_0/capacitors_1_6/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# VSUBS 2.34f
C99 cp1_buffer1_reverse_0/charge_pump1_reverse_0/capacitors_1_6/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# VSUBS 9.98f
C100 cp1_buffer1_reverse_0/charge_pump1_reverse_0/capacitors_1_6/capacitor_8_0/capacitor_7_0/buffer_digital_0/in VSUBS 2.61f
C101 cp1_buffer1_reverse_0/charge_pump1_reverse_0/capacitors_1_5/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# VSUBS 2.34f
C102 cp1_buffer1_reverse_0/charge_pump1_reverse_0/capacitors_1_5/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# VSUBS 9.98f
C103 cp1_buffer1_reverse_0/charge_pump1_reverse_0/capacitors_1_5/capacitor_8_0/capacitor_7_0/buffer_digital_0/in VSUBS 2.61f
C104 cp1_buffer1_reverse_0/charge_pump1_reverse_0/capacitors_1_4/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# VSUBS 2.34f
C105 cp1_buffer1_reverse_0/charge_pump1_reverse_0/capacitors_1_4/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# VSUBS 9.98f
C106 cp1_buffer1_reverse_0/charge_pump1_reverse_0/capacitors_1_4/capacitor_8_0/capacitor_7_0/buffer_digital_0/in VSUBS 2.61f
C107 cp1_buffer1_reverse_0/charge_pump1_reverse_0/capacitors_1_3/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# VSUBS 2.34f
C108 cp1_buffer1_reverse_0/charge_pump1_reverse_0/capacitors_1_3/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# VSUBS 9.98f
C109 cp1_buffer1_reverse_0/charge_pump1_reverse_0/capacitors_1_3/capacitor_8_0/capacitor_7_0/buffer_digital_0/in VSUBS 2.61f
C110 cp1_buffer1_2/charge_pump1_0/in6 VSUBS 11.4f
C111 cp1_buffer1_reverse_0/charge_pump1_reverse_0/capacitors_1_2/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# VSUBS 2.34f
C112 cp1_buffer1_reverse_0/charge_pump1_reverse_0/capacitors_1_2/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# VSUBS 9.98f
C113 cp1_buffer1_reverse_0/charge_pump1_reverse_0/capacitors_1_2/capacitor_8_0/capacitor_7_0/buffer_digital_0/in VSUBS 2.61f
C114 cp1_buffer1_reverse_0/charge_pump1_reverse_0/capacitors_1_1/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# VSUBS 2.34f
C115 cp1_buffer1_reverse_0/charge_pump1_reverse_0/capacitors_1_1/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# VSUBS 9.98f
C116 cp1_buffer1_reverse_0/charge_pump1_reverse_0/capacitors_1_1/capacitor_8_0/capacitor_7_0/buffer_digital_0/in VSUBS 2.61f
C117 cp1_buffer1_reverse_0/charge_pump1_reverse_0/capacitors_1_0/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# VSUBS 2.34f
C118 cp1_buffer1_reverse_0/charge_pump1_reverse_0/capacitors_1_0/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# VSUBS 9.98f
C119 cp1_buffer1_reverse_0/charge_pump1_reverse_0/capacitors_1_0/capacitor_8_0/capacitor_7_0/buffer_digital_0/in VSUBS 2.61f
C120 cp1_buffer1_reverse_0/charge_pump1_reverse_0/capacitor_8_1/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# VSUBS 2.34f
C121 cp1_buffer1_reverse_0/charge_pump1_reverse_0/clock_1/clk VSUBS 94.7f
C122 cp1_buffer1_reverse_0/charge_pump1_reverse_0/capacitor_8_1/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# VSUBS 9.98f
C123 cp1_buffer1_reverse_0/charge_pump1_reverse_0/capacitor_8_1/capacitor_7_0/buffer_digital_0/in VSUBS 2.61f
C124 cp1_buffer1_reverse_0/charge_pump1_reverse_0/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# VSUBS 2.34f
C125 cp1_buffer1_reverse_0/charge_pump1_reverse_0/clock_1/clkb VSUBS 0.101p
C126 cp1_buffer1_reverse_0/charge_pump1_reverse_0/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# VSUBS 9.98f
C127 cp1_buffer1_reverse_0/charge_pump1_reverse_0/capacitor_8_0/capacitor_7_0/buffer_digital_0/in VSUBS 2.61f
C128 cp1_buffer1_reverse_0/charge_pump1_reverse_0/clock_1/a_2432_n962# VSUBS 8.68f **FLOATING
C129 cp1_buffer1_reverse_0/charge_pump1_reverse_0/clock_1/a_2020_n482# VSUBS 2.57f **FLOATING
C130 cp1_buffer1_reverse_0/charge_pump1_reverse_0/clock_1/a_344_102# VSUBS 2.81f
C131 cp1_buffer1_reverse_0/charge_pump1_reverse_0/clock_1/a_2402_572# VSUBS 2.17f
C132 cp1_buffer1_reverse_0/charge_pump1_reverse_0/clock_1/a_344_n986# VSUBS 2.38f
C133 cp1_buffer1_1/clk_in VSUBS 6.57f
C134 cp1_buffer1_reverse_0/charge_pump1_reverse_0/clock_1/a_3246_118# VSUBS 6.83f
C135 cp1_buffer1_2/clk_out VSUBS 3.53f
C136 cp1_buffer1_2/charge_pump1_0/input1 VSUBS 22.5f
C137 cp1_buffer1_2/charge_pump1_0/input2 VSUBS 22.2f
C138 cp1_buffer1_2/charge_pump1_0/capacitors_1_12/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# VSUBS 2.34f
C139 cp1_buffer1_2/charge_pump1_0/capacitors_1_12/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# VSUBS 9.98f
C140 cp1_buffer1_2/charge_pump1_0/capacitors_1_12/capacitor_8_0/capacitor_7_0/buffer_digital_0/in VSUBS 2.61f
C141 cp1_buffer1_2/charge_pump1_0/capacitors_1_13/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# VSUBS 2.34f
C142 cp1_buffer1_2/charge_pump1_0/capacitors_1_13/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# VSUBS 9.98f
C143 cp1_buffer1_2/charge_pump1_0/capacitors_1_13/capacitor_8_0/capacitor_7_0/buffer_digital_0/in VSUBS 2.61f
C144 cp1_buffer1_2/charge_pump1_0/in4 VSUBS 11.4f
C145 cp1_buffer1_2/charge_pump1_0/capacitors_1_11/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# VSUBS 2.34f
C146 cp1_buffer1_2/charge_pump1_0/capacitors_1_11/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# VSUBS 9.98f
C147 cp1_buffer1_2/charge_pump1_0/capacitors_1_11/capacitor_8_0/capacitor_7_0/buffer_digital_0/in VSUBS 2.61f
C148 cp1_buffer1_2/charge_pump1_0/capacitors_1_10/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# VSUBS 2.34f
C149 cp1_buffer1_2/charge_pump1_0/capacitors_1_10/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# VSUBS 9.98f
C150 cp1_buffer1_2/charge_pump1_0/capacitors_1_10/capacitor_8_0/capacitor_7_0/buffer_digital_0/in VSUBS 2.61f
C151 cp1_buffer1_2/charge_pump1_0/m1_4341_n519# VSUBS 3.77f
C152 cp1_buffer1_2/charge_pump1_0/m1_12659_300# VSUBS 2.54f
C153 cp1_buffer1_2/charge_pump1_0/m1_12464_n576# VSUBS 4.26f
C154 cp1_buffer1_2/charge_pump1_0/capacitors_1_9/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# VSUBS 2.34f
C155 cp1_buffer1_2/charge_pump1_0/capacitors_1_9/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# VSUBS 9.98f
C156 cp1_buffer1_2/charge_pump1_0/capacitors_1_9/capacitor_8_0/capacitor_7_0/buffer_digital_0/in VSUBS 2.61f
C157 cp1_buffer1_2/charge_pump1_0/capacitors_1_8/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# VSUBS 2.34f
C158 cp1_buffer1_2/charge_pump1_0/capacitors_1_8/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# VSUBS 9.98f
C159 cp1_buffer1_2/charge_pump1_0/capacitors_1_8/capacitor_8_0/capacitor_7_0/buffer_digital_0/in VSUBS 2.61f
C160 cp1_buffer1_2/charge_pump1_0/capacitors_1_7/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# VSUBS 2.34f
C161 cp1_buffer1_2/charge_pump1_0/capacitors_1_7/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# VSUBS 9.98f
C162 cp1_buffer1_2/charge_pump1_0/capacitors_1_7/capacitor_8_0/capacitor_7_0/buffer_digital_0/in VSUBS 2.61f
C163 cp1_buffer1_2/charge_pump1_0/capacitors_1_6/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# VSUBS 2.34f
C164 cp1_buffer1_2/charge_pump1_0/capacitors_1_6/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# VSUBS 9.98f
C165 cp1_buffer1_2/charge_pump1_0/capacitors_1_6/capacitor_8_0/capacitor_7_0/buffer_digital_0/in VSUBS 2.61f
C166 cp1_buffer1_2/charge_pump1_0/capacitors_1_5/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# VSUBS 2.34f
C167 cp1_buffer1_2/charge_pump1_0/capacitors_1_5/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# VSUBS 9.98f
C168 cp1_buffer1_2/charge_pump1_0/capacitors_1_5/capacitor_8_0/capacitor_7_0/buffer_digital_0/in VSUBS 2.61f
C169 cp1_buffer1_2/charge_pump1_0/capacitors_1_4/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# VSUBS 2.34f
C170 cp1_buffer1_2/charge_pump1_0/capacitors_1_4/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# VSUBS 9.98f
C171 cp1_buffer1_2/charge_pump1_0/capacitors_1_4/capacitor_8_0/capacitor_7_0/buffer_digital_0/in VSUBS 2.61f
C172 cp1_buffer1_2/charge_pump1_0/capacitors_1_3/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# VSUBS 2.34f
C173 cp1_buffer1_2/charge_pump1_0/capacitors_1_3/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# VSUBS 9.98f
C174 cp1_buffer1_2/charge_pump1_0/capacitors_1_3/capacitor_8_0/capacitor_7_0/buffer_digital_0/in VSUBS 2.61f
C175 cp1_buffer1_2/charge_pump1_0/capacitors_1_2/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# VSUBS 2.34f
C176 cp1_buffer1_2/charge_pump1_0/capacitors_1_2/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# VSUBS 9.98f
C177 cp1_buffer1_2/charge_pump1_0/capacitors_1_2/capacitor_8_0/capacitor_7_0/buffer_digital_0/in VSUBS 2.61f
C178 cp1_buffer1_2/charge_pump1_0/capacitors_1_1/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# VSUBS 2.34f
C179 cp1_buffer1_2/charge_pump1_0/capacitors_1_1/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# VSUBS 9.98f
C180 cp1_buffer1_2/charge_pump1_0/capacitors_1_1/capacitor_8_0/capacitor_7_0/buffer_digital_0/in VSUBS 2.61f
C181 cp1_buffer1_2/charge_pump1_0/in1 VSUBS 10.9f
C182 cp1_buffer1_2/charge_pump1_0/capacitors_1_0/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# VSUBS 2.34f
C183 cp1_buffer1_2/charge_pump1_0/capacitors_1_0/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# VSUBS 9.98f
C184 cp1_buffer1_2/charge_pump1_0/capacitors_1_0/capacitor_8_0/capacitor_7_0/buffer_digital_0/in VSUBS 2.61f
C185 cp1_buffer1_2/charge_pump1_0/capacitor_8_1/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# VSUBS 2.34f
C186 cp1_buffer1_2/charge_pump1_0/clkb VSUBS 89.7f
C187 cp1_buffer1_2/charge_pump1_0/capacitor_8_1/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# VSUBS 9.98f
C188 cp1_buffer1_2/charge_pump1_0/capacitor_8_1/capacitor_7_0/buffer_digital_0/in VSUBS 2.61f
C189 cp1_buffer1_2/charge_pump1_0/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# VSUBS 2.34f
C190 cp1_buffer1_2/charge_pump1_0/clk VSUBS 89f
C191 cp1_buffer1_2/charge_pump1_0/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# VSUBS 9.98f
C192 cp1_buffer1_2/charge_pump1_0/capacitor_8_0/capacitor_7_0/buffer_digital_0/in VSUBS 2.61f
C193 cp1_buffer1_2/charge_pump1_0/clock_0/a_2432_n962# VSUBS 8.68f **FLOATING
C194 cp1_buffer1_2/charge_pump1_0/clock_0/a_2020_n482# VSUBS 2.57f **FLOATING
C195 cp1_buffer1_2/charge_pump1_0/clock_0/a_344_102# VSUBS 2.81f
C196 cp1_buffer1_2/charge_pump1_0/clock_0/a_2402_572# VSUBS 2.17f
C197 cp1_buffer1_2/charge_pump1_0/clock_0/a_344_n986# VSUBS 2.38f
C198 cp1_buffer1_2/charge_pump1_0/clock_0/a_3246_118# VSUBS 6.83f
C199 cp1_buffer1_2/charge_pump1_0/g2 VSUBS 2.34f
C200 cp1_buffer1_2/charge_pump1_0/vin VSUBS 13.4f
C201 cp1_buffer1_1/clk_out VSUBS 10.8f
C202 cp1_buffer1_1/charge_pump1_0/input1 VSUBS 22.5f
C203 cp1_buffer1_1/charge_pump1_0/input2 VSUBS 22.2f
C204 cp1_buffer1_1/charge_pump1_0/capacitors_1_12/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# VSUBS 2.34f
C205 cp1_buffer1_1/charge_pump1_0/capacitors_1_12/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# VSUBS 9.98f
C206 cp1_buffer1_1/charge_pump1_0/capacitors_1_12/capacitor_8_0/capacitor_7_0/buffer_digital_0/in VSUBS 2.61f
C207 cp1_buffer1_1/charge_pump1_0/capacitors_1_13/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# VSUBS 2.34f
C208 cp1_buffer1_1/charge_pump1_0/capacitors_1_13/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# VSUBS 9.98f
C209 cp1_buffer1_1/charge_pump1_0/capacitors_1_13/capacitor_8_0/capacitor_7_0/buffer_digital_0/in VSUBS 2.61f
C210 cp1_buffer1_1/charge_pump1_0/capacitors_1_11/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# VSUBS 2.34f
C211 cp1_buffer1_1/charge_pump1_0/capacitors_1_11/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# VSUBS 9.98f
C212 cp1_buffer1_1/charge_pump1_0/capacitors_1_11/capacitor_8_0/capacitor_7_0/buffer_digital_0/in VSUBS 2.61f
C213 cp1_buffer1_1/charge_pump1_0/capacitors_1_10/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# VSUBS 2.34f
C214 cp1_buffer1_1/charge_pump1_0/capacitors_1_10/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# VSUBS 9.98f
C215 cp1_buffer1_1/charge_pump1_0/capacitors_1_10/capacitor_8_0/capacitor_7_0/buffer_digital_0/in VSUBS 2.61f
C216 cp1_buffer1_1/charge_pump1_0/m1_4341_n519# VSUBS 3.77f
C217 cp1_buffer1_1/charge_pump1_0/m1_12659_300# VSUBS 2.54f
C218 cp1_buffer1_reverse_1/charge_pump1_reverse_0/nmos_dnw3_0/vs VSUBS 14.5f
C219 cp1_buffer1_1/charge_pump1_0/capacitors_1_9/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# VSUBS 2.34f
C220 cp1_buffer1_1/charge_pump1_0/capacitors_1_9/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# VSUBS 9.98f
C221 cp1_buffer1_1/charge_pump1_0/capacitors_1_9/capacitor_8_0/capacitor_7_0/buffer_digital_0/in VSUBS 2.61f
C222 cp1_buffer1_2/charge_pump1_0/in7 VSUBS 10.9f
C223 cp1_buffer1_1/charge_pump1_0/capacitors_1_8/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# VSUBS 2.34f
C224 cp1_buffer1_1/charge_pump1_0/capacitors_1_8/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# VSUBS 9.98f
C225 cp1_buffer1_1/charge_pump1_0/capacitors_1_8/capacitor_8_0/capacitor_7_0/buffer_digital_0/in VSUBS 2.61f
C226 cp1_buffer1_1/charge_pump1_0/capacitors_1_7/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# VSUBS 2.34f
C227 cp1_buffer1_1/charge_pump1_0/capacitors_1_7/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# VSUBS 9.98f
C228 cp1_buffer1_1/charge_pump1_0/capacitors_1_7/capacitor_8_0/capacitor_7_0/buffer_digital_0/in VSUBS 2.61f
C229 cp1_buffer1_1/charge_pump1_0/capacitors_1_6/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# VSUBS 2.34f
C230 cp1_buffer1_1/charge_pump1_0/capacitors_1_6/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# VSUBS 9.98f
C231 cp1_buffer1_1/charge_pump1_0/capacitors_1_6/capacitor_8_0/capacitor_7_0/buffer_digital_0/in VSUBS 2.61f
C232 cp1_buffer1_1/charge_pump1_0/capacitors_1_5/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# VSUBS 2.34f
C233 cp1_buffer1_1/charge_pump1_0/capacitors_1_5/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# VSUBS 9.98f
C234 cp1_buffer1_1/charge_pump1_0/capacitors_1_5/capacitor_8_0/capacitor_7_0/buffer_digital_0/in VSUBS 2.61f
C235 cp1_buffer1_1/charge_pump1_0/capacitors_1_4/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# VSUBS 2.34f
C236 cp1_buffer1_1/charge_pump1_0/capacitors_1_4/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# VSUBS 9.98f
C237 cp1_buffer1_1/charge_pump1_0/capacitors_1_4/capacitor_8_0/capacitor_7_0/buffer_digital_0/in VSUBS 2.61f
C238 cp1_buffer1_2/charge_pump1_0/in2 VSUBS 11.3f
C239 cp1_buffer1_1/charge_pump1_0/capacitors_1_3/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# VSUBS 2.34f
C240 cp1_buffer1_1/charge_pump1_0/capacitors_1_3/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# VSUBS 9.98f
C241 cp1_buffer1_1/charge_pump1_0/capacitors_1_3/capacitor_8_0/capacitor_7_0/buffer_digital_0/in VSUBS 2.61f
C242 cp1_buffer1_2/charge_pump1_0/in3 VSUBS 11.2f
C243 cp1_buffer1_1/charge_pump1_0/capacitors_1_2/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# VSUBS 2.34f
C244 cp1_buffer1_1/charge_pump1_0/capacitors_1_2/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# VSUBS 9.98f
C245 cp1_buffer1_1/charge_pump1_0/capacitors_1_2/capacitor_8_0/capacitor_7_0/buffer_digital_0/in VSUBS 2.61f
C246 cp1_buffer1_1/charge_pump1_0/capacitors_1_1/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# VSUBS 2.34f
C247 cp1_buffer1_1/charge_pump1_0/capacitors_1_1/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# VSUBS 9.98f
C248 cp1_buffer1_1/charge_pump1_0/capacitors_1_1/capacitor_8_0/capacitor_7_0/buffer_digital_0/in VSUBS 2.61f
C249 cp1_buffer1_1/charge_pump1_0/capacitors_1_0/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# VSUBS 2.34f
C250 cp1_buffer1_1/charge_pump1_0/capacitors_1_0/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# VSUBS 9.98f
C251 cp1_buffer1_1/charge_pump1_0/capacitors_1_0/capacitor_8_0/capacitor_7_0/buffer_digital_0/in VSUBS 2.61f
C252 cp1_buffer1_1/charge_pump1_0/capacitor_8_1/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# VSUBS 2.34f
C253 cp1_buffer1_1/charge_pump1_0/clkb VSUBS 89.8f
C254 cp1_buffer1_1/charge_pump1_0/capacitor_8_1/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# VSUBS 9.98f
C255 cp1_buffer1_1/charge_pump1_0/capacitor_8_1/capacitor_7_0/buffer_digital_0/in VSUBS 2.61f
C256 cp1_buffer1_1/charge_pump1_0/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# VSUBS 2.34f
C257 cp1_buffer1_1/charge_pump1_0/clk VSUBS 89.1f
C258 cp1_buffer1_1/charge_pump1_0/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# VSUBS 9.98f
C259 cp1_buffer1_1/charge_pump1_0/capacitor_8_0/capacitor_7_0/buffer_digital_0/in VSUBS 2.61f
C260 cp1_buffer1_1/charge_pump1_0/clock_0/a_2432_n962# VSUBS 8.68f **FLOATING
C261 cp1_buffer1_1/charge_pump1_0/clock_0/a_2020_n482# VSUBS 2.57f **FLOATING
C262 cp1_buffer1_1/charge_pump1_0/clock_0/a_344_102# VSUBS 2.81f
C263 cp1_buffer1_1/charge_pump1_0/clock_0/a_2402_572# VSUBS 2.17f
C264 cp1_buffer1_1/charge_pump1_0/clock_0/a_344_n986# VSUBS 2.38f
C265 cp1_buffer1_1/charge_pump1_0/clock_0/a_3246_118# VSUBS 6.83f
C266 cp1_buffer1_1/charge_pump1_0/g2 VSUBS 2.34f
C267 cp1_buffer1_1/charge_pump1_0/vin VSUBS 13.3f
C268 cp1_buffer1_0/clk_in VSUBS 2.92f
C269 cp1_buffer1_0/clk_out VSUBS 10.6f
C270 cp1_buffer1_0/charge_pump1_0/input1 VSUBS 22.5f
C271 cp1_buffer1_0/charge_pump1_0/input2 VSUBS 22.2f
C272 cp1_buffer1_0/charge_pump1_0/capacitors_1_12/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# VSUBS 2.34f
C273 cp1_buffer1_0/charge_pump1_0/capacitors_1_12/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# VSUBS 9.98f
C274 cp1_buffer1_0/charge_pump1_0/capacitors_1_12/capacitor_8_0/capacitor_7_0/buffer_digital_0/in VSUBS 2.61f
C275 cp1_buffer1_2/charge_pump1_0/in5 VSUBS 11.3f
C276 cp1_buffer1_0/charge_pump1_0/capacitors_1_13/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# VSUBS 2.34f
C277 cp1_buffer1_0/charge_pump1_0/capacitors_1_13/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# VSUBS 9.98f
C278 cp1_buffer1_0/charge_pump1_0/capacitors_1_13/capacitor_8_0/capacitor_7_0/buffer_digital_0/in VSUBS 2.61f
C279 cp1_buffer1_0/charge_pump1_0/capacitors_1_11/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# VSUBS 2.34f
C280 cp1_buffer1_0/charge_pump1_0/capacitors_1_11/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# VSUBS 9.98f
C281 cp1_buffer1_0/charge_pump1_0/capacitors_1_11/capacitor_8_0/capacitor_7_0/buffer_digital_0/in VSUBS 2.61f
C282 cp1_buffer1_0/charge_pump1_0/capacitors_1_10/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# VSUBS 2.34f
C283 cp1_buffer1_0/charge_pump1_0/capacitors_1_10/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# VSUBS 9.98f
C284 cp1_buffer1_0/charge_pump1_0/capacitors_1_10/capacitor_8_0/capacitor_7_0/buffer_digital_0/in VSUBS 2.61f
C285 cp1_buffer1_0/charge_pump1_0/m1_4341_n519# VSUBS 3.77f
C286 cp1_buffer1_0/charge_pump1_0/m1_12659_300# VSUBS 2.54f
C287 cp1_buffer1_reverse_0/charge_pump1_reverse_0/nmos_dnw3_0/vs VSUBS 14.7f
C288 cp1_buffer1_0/charge_pump1_0/capacitors_1_9/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# VSUBS 2.34f
C289 cp1_buffer1_0/charge_pump1_0/capacitors_1_9/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# VSUBS 9.99f
C290 cp1_buffer1_0/charge_pump1_0/capacitors_1_9/capacitor_8_0/capacitor_7_0/buffer_digital_0/in VSUBS 2.61f
C291 cp1_buffer1_0/charge_pump1_0/capacitors_1_8/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# VSUBS 2.34f
C292 cp1_buffer1_0/charge_pump1_0/capacitors_1_8/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# VSUBS 9.98f
C293 cp1_buffer1_0/charge_pump1_0/capacitors_1_8/capacitor_8_0/capacitor_7_0/buffer_digital_0/in VSUBS 2.61f
C294 cp1_buffer1_0/charge_pump1_0/capacitors_1_7/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# VSUBS 2.34f
C295 cp1_buffer1_0/charge_pump1_0/capacitors_1_7/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# VSUBS 9.98f
C296 cp1_buffer1_0/charge_pump1_0/capacitors_1_7/capacitor_8_0/capacitor_7_0/buffer_digital_0/in VSUBS 2.61f
C297 cp1_buffer1_0/charge_pump1_0/capacitors_1_6/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# VSUBS 2.34f
C298 cp1_buffer1_0/charge_pump1_0/capacitors_1_6/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# VSUBS 9.98f
C299 cp1_buffer1_0/charge_pump1_0/capacitors_1_6/capacitor_8_0/capacitor_7_0/buffer_digital_0/in VSUBS 2.61f
C300 cp1_buffer1_0/charge_pump1_0/capacitors_1_5/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# VSUBS 2.34f
C301 cp1_buffer1_0/charge_pump1_0/capacitors_1_5/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# VSUBS 9.98f
C302 cp1_buffer1_0/charge_pump1_0/capacitors_1_5/capacitor_8_0/capacitor_7_0/buffer_digital_0/in VSUBS 2.61f
C303 cp1_buffer1_0/charge_pump1_0/capacitors_1_4/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# VSUBS 2.34f
C304 cp1_buffer1_0/charge_pump1_0/capacitors_1_4/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# VSUBS 9.98f
C305 cp1_buffer1_0/charge_pump1_0/capacitors_1_4/capacitor_8_0/capacitor_7_0/buffer_digital_0/in VSUBS 2.61f
C306 cp1_buffer1_0/charge_pump1_0/capacitors_1_3/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# VSUBS 2.34f
C307 cp1_buffer1_0/charge_pump1_0/capacitors_1_3/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# VSUBS 9.98f
C308 cp1_buffer1_0/charge_pump1_0/capacitors_1_3/capacitor_8_0/capacitor_7_0/buffer_digital_0/in VSUBS 2.61f
C309 cp1_buffer1_0/charge_pump1_0/capacitors_1_2/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# VSUBS 2.34f
C310 cp1_buffer1_0/charge_pump1_0/capacitors_1_2/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# VSUBS 9.98f
C311 cp1_buffer1_0/charge_pump1_0/capacitors_1_2/capacitor_8_0/capacitor_7_0/buffer_digital_0/in VSUBS 2.61f
C312 cp1_buffer1_0/charge_pump1_0/capacitors_1_1/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# VSUBS 2.34f
C313 cp1_buffer1_0/charge_pump1_0/capacitors_1_1/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# VSUBS 9.98f
C314 cp1_buffer1_0/charge_pump1_0/capacitors_1_1/capacitor_8_0/capacitor_7_0/buffer_digital_0/in VSUBS 2.61f
C315 cp1_buffer1_0/charge_pump1_0/capacitors_1_0/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# VSUBS 2.34f
C316 cp1_buffer1_0/charge_pump1_0/capacitors_1_0/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# VSUBS 9.98f
C317 cp1_buffer1_0/charge_pump1_0/capacitors_1_0/capacitor_8_0/capacitor_7_0/buffer_digital_0/in VSUBS 2.61f
C318 cp1_buffer1_0/charge_pump1_0/capacitor_8_1/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# VSUBS 2.34f
C319 cp1_buffer1_0/charge_pump1_0/clkb VSUBS 89.8f
C320 cp1_buffer1_0/charge_pump1_0/capacitor_8_1/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# VSUBS 9.98f
C321 cp1_buffer1_0/charge_pump1_0/capacitor_8_1/capacitor_7_0/buffer_digital_0/in VSUBS 2.61f
C322 cp1_buffer1_0/charge_pump1_0/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# VSUBS 2.34f
C323 cp1_buffer1_0/charge_pump1_0/clk VSUBS 88.9f
C324 cp1_buffer1_2/vdd VSUBS 2.86p
C325 cp1_buffer1_0/charge_pump1_0/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# VSUBS 9.98f
C326 cp1_buffer1_0/charge_pump1_0/capacitor_8_0/capacitor_7_0/buffer_digital_0/in VSUBS 2.61f
C327 cp1_buffer1_0/charge_pump1_0/clock_0/a_2432_n962# VSUBS 8.68f **FLOATING
C328 cp1_buffer1_0/charge_pump1_0/clock_0/a_2020_n482# VSUBS 2.57f **FLOATING
C329 cp1_buffer1_0/charge_pump1_0/clock_0/a_344_102# VSUBS 2.81f
C330 cp1_buffer1_0/charge_pump1_0/clock_0/a_2402_572# VSUBS 2.17f
C331 cp1_buffer1_0/charge_pump1_0/clock_0/a_344_n986# VSUBS 2.38f
C332 cp1_buffer1_0/charge_pump1_0/clock_0/a_3246_118# VSUBS 6.83f
C333 cp1_buffer1_0/charge_pump1_0/g2 VSUBS 2.34f
C334 cp1_buffer1_0/charge_pump1_0/vin VSUBS 10.4f
.ends

.subckt sky130_fd_pr__nfet_01v8_D4CMYK a_15_n130# a_63_n42# a_n177_n130# a_255_n42#
+ a_n129_n42# a_111_64# a_n321_n42# a_159_n42# a_n81_64# a_n273_64# a_351_n42# a_207_n130#
+ a_303_64# a_n33_n42# a_n369_n130# a_n225_n42# a_n413_n42# VSUBS
X0 a_63_n42# a_15_n130# a_n33_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X1 a_n33_n42# a_n81_64# a_n129_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X2 a_351_n42# a_303_64# a_255_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X3 a_159_n42# a_111_64# a_63_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X4 a_255_n42# a_207_n130# a_159_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X5 a_n321_n42# a_n369_n130# a_n413_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X6 a_n225_n42# a_n273_64# a_n321_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X7 a_n129_n42# a_n177_n130# a_n225_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
.ends

.subckt capacitor_5 cp_clk i1 vd2 vd1 vd4 vd3 clk GND VDD
Xbuffer_digital_1 i1 buffer_digital_1/in VDD GND buffer_digital
Xsky130_fd_pr__nfet_01v8_D4CMYK_0 vd2 GND vd2 GND GND vd2 GND GND vd2 vd2 GND vd2
+ vd2 GND vd2 GND GND GND sky130_fd_pr__nfet_01v8_D4CMYK
Xsky130_fd_pr__pfet_01v8_4ZKXAA_1 vd3 vd3 GND vd3 vd3 GND vd3 GND vd3 GND GND vd3
+ GND vd3 vd3 GND GND vd3 vd3 GND vd3 GND GND sky130_fd_pr__pfet_01v8_4ZKXAA
Xsky130_fd_pr__pfet_01v8_4ZKXAA_2 vd4 vd4 GND vd4 vd4 GND vd4 GND vd4 GND GND vd4
+ GND vd4 vd4 GND GND vd4 vd4 GND vd4 GND GND sky130_fd_pr__pfet_01v8_4ZKXAA
Xsky130_fd_pr__pfet_01v8_4ZKXAA_3 vd3 vd3 GND vd3 vd3 GND vd3 GND vd3 GND GND vd3
+ GND vd3 vd3 GND GND vd3 vd3 GND vd3 GND GND sky130_fd_pr__pfet_01v8_4ZKXAA
Xsky130_fd_pr__nfet_01v8_NJGC45_0 GND vd1 GND vd1 vd1 GND GND vd1 vd1 GND vd1 GND
+ GND GND GND GND vd1 GND vd1 vd1 vd1 GND sky130_fd_pr__nfet_01v8_NJGC45
Xbuffer_and_gate_0 buffer_digital_1/in clk buffer_and_gate_0/out GND VDD buffer_and_gate
X0 buffer_and_gate_0/out cp_clk sky130_fd_pr__cap_mim_m3_1 l=4.97 w=5
C0 buffer_digital_1/in i1 2.94f
C1 buffer_and_gate_0/and_gate_0/a_n78_396# GND 2.36f
C2 clk GND 8.64f
C3 VDD GND 21f
C4 buffer_and_gate_0/buffer_0/a_1436_1552# GND 10.2f
C5 vd1 GND 3.43f
C6 vd3 GND 7.1f
C7 vd4 GND 2.86f
C8 vd2 GND 3.08f
C9 buffer_digital_1/in GND 2.67f
.ends

.subckt capacitors_5 capacitor_5_7/i1 capacitor_5_1/i1 capacitor_5_6/i1 capacitor_5_0/i1
+ capacitor_5_7/vd4 capacitor_5_3/i1 capacitor_5_7/vd2 capacitor_5_7/vd1 capacitor_5_7/cp_clk
+ capacitor_5_4/i1 capacitor_5_2/i1 capacitor_5_7/clk capacitor_5_7/vd3 capacitor_5_5/i1
+ VSUBS capacitor_5_7/VDD
Xcapacitor_5_5 capacitor_5_7/cp_clk capacitor_5_5/i1 capacitor_5_7/VDD capacitor_5_7/VDD
+ capacitor_5_7/VDD capacitor_5_7/VDD capacitor_5_7/clk VSUBS capacitor_5_7/VDD capacitor_5
Xcapacitor_5_6 capacitor_5_7/cp_clk capacitor_5_6/i1 capacitor_5_7/VDD capacitor_5_7/VDD
+ capacitor_5_7/VDD capacitor_5_7/VDD capacitor_5_7/clk VSUBS capacitor_5_7/VDD capacitor_5
Xcapacitor_5_7 capacitor_5_7/cp_clk capacitor_5_7/i1 capacitor_5_7/vd2 capacitor_5_7/vd1
+ capacitor_5_7/vd4 capacitor_5_7/vd3 capacitor_5_7/clk VSUBS capacitor_5_7/VDD capacitor_5
Xcapacitor_5_0 capacitor_5_7/cp_clk capacitor_5_0/i1 capacitor_5_7/VDD capacitor_5_7/VDD
+ capacitor_5_7/VDD capacitor_5_7/VDD capacitor_5_7/clk VSUBS capacitor_5_7/VDD capacitor_5
Xcapacitor_5_1 capacitor_5_7/cp_clk capacitor_5_1/i1 capacitor_5_7/VDD capacitor_5_7/VDD
+ capacitor_5_7/VDD capacitor_5_7/VDD capacitor_5_7/clk VSUBS capacitor_5_7/VDD capacitor_5
Xcapacitor_5_2 capacitor_5_7/cp_clk capacitor_5_2/i1 capacitor_5_7/VDD capacitor_5_7/VDD
+ capacitor_5_7/VDD capacitor_5_7/VDD capacitor_5_7/clk VSUBS capacitor_5_7/VDD capacitor_5
Xcapacitor_5_3 capacitor_5_7/cp_clk capacitor_5_3/i1 capacitor_5_7/VDD capacitor_5_7/VDD
+ capacitor_5_7/VDD capacitor_5_7/VDD capacitor_5_7/clk VSUBS capacitor_5_7/VDD capacitor_5
Xcapacitor_5_4 capacitor_5_7/cp_clk capacitor_5_4/i1 capacitor_5_7/VDD capacitor_5_7/VDD
+ capacitor_5_7/VDD capacitor_5_7/VDD capacitor_5_7/clk VSUBS capacitor_5_7/VDD capacitor_5
C0 capacitor_5_7/cp_clk capacitor_5_7/VDD 11.7f
C1 capacitor_5_7/clk capacitor_5_7/VDD 13f
C2 capacitor_5_4/buffer_and_gate_0/and_gate_0/a_n78_396# VSUBS 2.38f
C3 capacitor_5_4/buffer_and_gate_0/buffer_0/a_1436_1552# VSUBS 10.1f
C4 capacitor_5_4/buffer_digital_1/in VSUBS 2.64f
C5 capacitor_5_3/buffer_and_gate_0/and_gate_0/a_n78_396# VSUBS 2.37f
C6 capacitor_5_3/buffer_and_gate_0/buffer_0/a_1436_1552# VSUBS 10.1f
C7 capacitor_5_3/buffer_digital_1/in VSUBS 2.64f
C8 capacitor_5_2/buffer_and_gate_0/and_gate_0/a_n78_396# VSUBS 2.38f
C9 capacitor_5_2/buffer_and_gate_0/buffer_0/a_1436_1552# VSUBS 10.1f
C10 capacitor_5_2/buffer_digital_1/in VSUBS 2.64f
C11 capacitor_5_1/buffer_and_gate_0/and_gate_0/a_n78_396# VSUBS 2.38f
C12 capacitor_5_1/buffer_and_gate_0/buffer_0/a_1436_1552# VSUBS 10.1f
C13 capacitor_5_1/buffer_digital_1/in VSUBS 2.64f
C14 capacitor_5_0/buffer_and_gate_0/and_gate_0/a_n78_396# VSUBS 2.34f
C15 capacitor_5_0/buffer_and_gate_0/buffer_0/a_1436_1552# VSUBS 9.98f
C16 capacitor_5_0/buffer_digital_1/in VSUBS 2.58f
C17 capacitor_5_7/cp_clk VSUBS 20.1f
C18 capacitor_5_7/buffer_and_gate_0/and_gate_0/a_n78_396# VSUBS 2.38f
C19 capacitor_5_7/clk VSUBS 71.2f
C20 capacitor_5_7/VDD VSUBS 0.26p
C21 capacitor_5_7/buffer_and_gate_0/buffer_0/a_1436_1552# VSUBS 10.1f
C22 capacitor_5_7/vd1 VSUBS 2.32f
C23 capacitor_5_7/vd3 VSUBS 3.83f
C24 capacitor_5_7/vd2 VSUBS 2.22f
C25 capacitor_5_7/buffer_digital_1/in VSUBS 2.64f
C26 capacitor_5_6/buffer_and_gate_0/and_gate_0/a_n78_396# VSUBS 2.38f
C27 capacitor_5_6/buffer_and_gate_0/buffer_0/a_1436_1552# VSUBS 10.1f
C28 capacitor_5_6/buffer_digital_1/in VSUBS 2.64f
C29 capacitor_5_5/buffer_and_gate_0/and_gate_0/a_n78_396# VSUBS 2.38f
C30 capacitor_5_5/buffer_and_gate_0/buffer_0/a_1436_1552# VSUBS 10.1f
C31 capacitor_5_5/buffer_digital_1/in VSUBS 2.64f
.ends

.subckt nmos_diode2 a_350_n764# a_970_n762# a_410_n892# dw_118_n1078# VSUBS
X0 a_410_n892# a_410_n892# a_350_n764# dw_118_n1078# sky130_fd_pr__nfet_01v8 ad=0.873 pd=6.6 as=0.903 ps=6.62 w=3.01 l=1
X1 a_350_n764# a_970_n762# a_970_n762# dw_118_n1078# sky130_fd_pr__nfet_01v8 ad=0.993 pd=6.68 as=0.873 ps=6.6 w=3.01 l=1
C0 dw_118_n1078# VSUBS 8.16f
.ends

.subckt charge_pump in1 in3 in5 input1 input2 out clk clkb clk_in g1 g2 vin a_18057_18271#
+ in6 in8 in4 in7 in2 vs clock_0/gnd clock_0/vdd
Xsky130_fd_pr__cap_mim_m3_1_MH6KF8_4 g1 clk clock_0/gnd sky130_fd_pr__cap_mim_m3_1_MH6KF8
Xsky130_fd_pr__cap_mim_m3_1_MH6KF8_5 g2 clkb clock_0/gnd sky130_fd_pr__cap_mim_m3_1_MH6KF8
Xcapacitors_5_1 in8 in2 in7 in1 clock_0/vdd in4 clock_0/vdd clock_0/vdd input2 in5
+ in3 clkb clock_0/vdd in6 clock_0/gnd clock_0/vdd capacitors_5
Xcapacitors_5_0 in8 in2 in7 in1 clock_0/vdd in4 clock_0/vdd clock_0/vdd input1 in5
+ in3 clk clock_0/vdd in6 clock_0/gnd clock_0/vdd capacitors_5
Xnmos_dnw3_0 vin input1 input2 g1 g2 vs clock_0/gnd nmos_dnw3
Xclock_0 clk_in clock_0/vdd clock_0/gnd clk clkb clock
Xsky130_fd_pr__pfet_01v8_4RPJ49_0 clock_0/gnd clock_0/vdd clock_0/vdd clock_0/gnd
+ clock_0/gnd clock_0/vdd clock_0/vdd clock_0/vdd clock_0/gnd clock_0/vdd clock_0/gnd
+ clock_0/gnd clock_0/vdd clock_0/gnd clock_0/gnd clock_0/gnd clock_0/vdd clock_0/vdd
+ clock_0/vdd clock_0/vdd clock_0/gnd clock_0/vdd clock_0/gnd clock_0/gnd clock_0/gnd
+ clock_0/gnd clock_0/gnd clock_0/gnd clock_0/gnd clock_0/vdd clock_0/gnd clock_0/vdd
+ clock_0/gnd clock_0/gnd clock_0/vdd clock_0/gnd clock_0/gnd clock_0/vdd clock_0/vdd
+ clock_0/gnd clock_0/vdd clock_0/gnd clock_0/gnd clock_0/vdd clock_0/gnd clock_0/gnd
+ clock_0/vdd clock_0/vdd clock_0/gnd clock_0/gnd clock_0/vdd clock_0/vdd clock_0/vdd
+ clock_0/gnd clock_0/gnd clock_0/vdd clock_0/vdd clock_0/gnd clock_0/gnd clock_0/vdd
+ clock_0/vdd clock_0/gnd clock_0/vdd clock_0/gnd clock_0/vdd clock_0/gnd clock_0/gnd
+ clock_0/gnd clock_0/vdd clock_0/gnd clock_0/gnd clock_0/gnd clock_0/vdd clock_0/vdd
+ clock_0/gnd clock_0/gnd clock_0/vdd clock_0/vdd clock_0/gnd clock_0/gnd clock_0/vdd
+ clock_0/vdd clock_0/gnd clock_0/gnd clock_0/gnd clock_0/vdd clock_0/vdd clock_0/vdd
+ clock_0/vdd clock_0/vdd clock_0/vdd clock_0/vdd clock_0/vdd clock_0/vdd clock_0/gnd
+ clock_0/gnd clock_0/vdd clock_0/vdd clock_0/vdd clock_0/gnd clock_0/vdd clock_0/vdd
+ clock_0/vdd clock_0/vdd clock_0/vdd clock_0/gnd clock_0/vdd clock_0/vdd clock_0/gnd
+ clock_0/vdd clock_0/vdd clock_0/gnd clock_0/gnd clock_0/gnd clock_0/gnd clock_0/gnd
+ clock_0/vdd clock_0/vdd clock_0/vdd clock_0/gnd clock_0/vdd clock_0/vdd clock_0/gnd
+ clock_0/vdd clock_0/gnd clock_0/vdd clock_0/vdd clock_0/vdd clock_0/gnd clock_0/gnd
+ clock_0/vdd clock_0/vdd clock_0/gnd clock_0/vdd clock_0/vdd clock_0/vdd clock_0/vdd
+ clock_0/gnd clock_0/vdd clock_0/gnd clock_0/gnd clock_0/gnd clock_0/vdd clock_0/vdd
+ clock_0/vdd clock_0/gnd clock_0/gnd clock_0/gnd clock_0/gnd clock_0/vdd clock_0/gnd
+ clock_0/gnd clock_0/gnd clock_0/vdd clock_0/gnd clock_0/gnd clock_0/gnd clock_0/gnd
+ clock_0/vdd clock_0/gnd clock_0/gnd clock_0/vdd clock_0/vdd sky130_fd_pr__pfet_01v8_4RPJ49
Xsky130_fd_pr__pfet_01v8_4RPJ49_1 clock_0/gnd clock_0/vdd clock_0/vdd clock_0/gnd
+ clock_0/gnd clock_0/vdd clock_0/vdd clock_0/vdd clock_0/gnd clock_0/vdd clock_0/gnd
+ clock_0/gnd clock_0/vdd clock_0/gnd clock_0/gnd clock_0/gnd clock_0/vdd clock_0/vdd
+ clock_0/vdd clock_0/vdd clock_0/gnd clock_0/vdd clock_0/gnd clock_0/gnd clock_0/gnd
+ clock_0/gnd clock_0/gnd clock_0/gnd clock_0/gnd clock_0/vdd clock_0/gnd clock_0/vdd
+ clock_0/gnd clock_0/gnd clock_0/vdd clock_0/gnd clock_0/gnd clock_0/vdd clock_0/vdd
+ clock_0/gnd clock_0/vdd clock_0/gnd clock_0/gnd clock_0/vdd clock_0/gnd clock_0/gnd
+ clock_0/vdd clock_0/vdd clock_0/gnd clock_0/gnd clock_0/vdd clock_0/vdd clock_0/vdd
+ clock_0/gnd clock_0/gnd clock_0/vdd clock_0/vdd clock_0/gnd clock_0/gnd clock_0/vdd
+ clock_0/vdd clock_0/gnd clock_0/vdd clock_0/gnd clock_0/vdd clock_0/gnd clock_0/gnd
+ clock_0/gnd clock_0/vdd clock_0/gnd clock_0/gnd clock_0/gnd clock_0/vdd clock_0/vdd
+ clock_0/gnd clock_0/gnd clock_0/vdd clock_0/vdd clock_0/gnd clock_0/gnd clock_0/vdd
+ clock_0/vdd clock_0/gnd clock_0/gnd clock_0/gnd clock_0/vdd clock_0/vdd clock_0/vdd
+ clock_0/vdd clock_0/vdd clock_0/vdd clock_0/vdd clock_0/vdd clock_0/vdd clock_0/gnd
+ clock_0/gnd clock_0/vdd clock_0/vdd clock_0/vdd clock_0/gnd clock_0/vdd clock_0/vdd
+ clock_0/vdd clock_0/vdd clock_0/vdd clock_0/gnd clock_0/vdd clock_0/vdd clock_0/gnd
+ clock_0/vdd clock_0/vdd clock_0/gnd clock_0/gnd clock_0/gnd clock_0/gnd clock_0/gnd
+ clock_0/vdd clock_0/vdd clock_0/vdd clock_0/gnd clock_0/vdd clock_0/vdd clock_0/gnd
+ clock_0/vdd clock_0/gnd clock_0/vdd clock_0/vdd clock_0/vdd clock_0/gnd clock_0/gnd
+ clock_0/vdd clock_0/vdd clock_0/gnd clock_0/vdd clock_0/vdd clock_0/vdd clock_0/vdd
+ clock_0/gnd clock_0/vdd clock_0/gnd clock_0/gnd clock_0/gnd clock_0/vdd clock_0/vdd
+ clock_0/vdd clock_0/gnd clock_0/gnd clock_0/gnd clock_0/gnd clock_0/vdd clock_0/gnd
+ clock_0/gnd clock_0/gnd clock_0/vdd clock_0/gnd clock_0/gnd clock_0/gnd clock_0/gnd
+ clock_0/vdd clock_0/gnd clock_0/gnd clock_0/vdd clock_0/vdd sky130_fd_pr__pfet_01v8_4RPJ49
Xsky130_fd_pr__nfet_01v8_NJGC8F_0 clock_0/vdd clock_0/gnd clock_0/gnd clock_0/vdd
+ clock_0/vdd clock_0/gnd clock_0/gnd clock_0/vdd clock_0/gnd clock_0/vdd clock_0/gnd
+ clock_0/gnd clock_0/vdd clock_0/gnd clock_0/gnd clock_0/gnd clock_0/vdd clock_0/gnd
+ clock_0/vdd clock_0/vdd clock_0/gnd clock_0/vdd clock_0/vdd clock_0/vdd clock_0/vdd
+ clock_0/gnd clock_0/vdd clock_0/vdd clock_0/gnd clock_0/vdd clock_0/vdd clock_0/gnd
+ clock_0/gnd clock_0/gnd clock_0/gnd clock_0/gnd clock_0/vdd clock_0/gnd clock_0/gnd
+ clock_0/vdd clock_0/gnd clock_0/gnd clock_0/gnd clock_0/vdd clock_0/gnd clock_0/gnd
+ clock_0/vdd clock_0/gnd clock_0/gnd clock_0/gnd clock_0/vdd clock_0/vdd clock_0/gnd
+ clock_0/gnd clock_0/vdd clock_0/gnd clock_0/gnd clock_0/vdd clock_0/gnd clock_0/gnd
+ clock_0/gnd clock_0/vdd clock_0/vdd clock_0/vdd clock_0/gnd clock_0/gnd clock_0/gnd
+ clock_0/gnd clock_0/vdd clock_0/gnd clock_0/vdd clock_0/gnd clock_0/vdd clock_0/gnd
+ clock_0/gnd clock_0/vdd clock_0/gnd clock_0/vdd clock_0/vdd clock_0/vdd clock_0/vdd
+ clock_0/vdd clock_0/vdd clock_0/gnd clock_0/gnd clock_0/gnd clock_0/gnd clock_0/gnd
+ clock_0/vdd clock_0/gnd clock_0/gnd clock_0/vdd clock_0/vdd clock_0/gnd clock_0/vdd
+ clock_0/vdd clock_0/vdd clock_0/vdd clock_0/gnd clock_0/vdd clock_0/gnd clock_0/gnd
+ clock_0/gnd clock_0/gnd clock_0/gnd clock_0/vdd clock_0/vdd clock_0/vdd clock_0/vdd
+ clock_0/gnd clock_0/vdd clock_0/vdd clock_0/vdd clock_0/vdd clock_0/gnd clock_0/vdd
+ clock_0/gnd clock_0/vdd clock_0/vdd clock_0/gnd clock_0/gnd clock_0/vdd clock_0/gnd
+ clock_0/gnd clock_0/vdd clock_0/vdd clock_0/vdd clock_0/gnd clock_0/gnd clock_0/vdd
+ clock_0/gnd clock_0/gnd clock_0/gnd clock_0/vdd clock_0/vdd clock_0/gnd clock_0/vdd
+ clock_0/vdd clock_0/vdd clock_0/gnd clock_0/vdd clock_0/vdd clock_0/gnd clock_0/gnd
+ clock_0/gnd clock_0/vdd clock_0/vdd clock_0/vdd clock_0/gnd clock_0/vdd clock_0/vdd
+ clock_0/vdd clock_0/vdd clock_0/vdd clock_0/vdd clock_0/gnd clock_0/vdd clock_0/gnd
+ clock_0/vdd clock_0/gnd clock_0/gnd clock_0/gnd sky130_fd_pr__nfet_01v8_NJGC8F
Xsky130_fd_pr__nfet_01v8_NJGC8F_1 clock_0/vdd clock_0/gnd clock_0/gnd clock_0/vdd
+ clock_0/vdd clock_0/gnd clock_0/gnd clock_0/vdd clock_0/gnd clock_0/vdd clock_0/gnd
+ clock_0/gnd clock_0/vdd clock_0/gnd clock_0/gnd clock_0/gnd clock_0/vdd clock_0/gnd
+ clock_0/vdd clock_0/vdd clock_0/gnd clock_0/vdd clock_0/vdd clock_0/vdd clock_0/vdd
+ clock_0/gnd clock_0/vdd clock_0/vdd clock_0/gnd clock_0/vdd clock_0/vdd clock_0/gnd
+ clock_0/gnd clock_0/gnd clock_0/gnd clock_0/gnd clock_0/vdd clock_0/gnd clock_0/gnd
+ clock_0/vdd clock_0/gnd clock_0/gnd clock_0/gnd clock_0/vdd clock_0/gnd clock_0/gnd
+ clock_0/vdd clock_0/gnd clock_0/gnd clock_0/gnd clock_0/vdd clock_0/vdd clock_0/gnd
+ clock_0/gnd clock_0/vdd clock_0/gnd clock_0/gnd clock_0/vdd clock_0/gnd clock_0/gnd
+ clock_0/gnd clock_0/vdd clock_0/vdd clock_0/vdd clock_0/gnd clock_0/gnd clock_0/gnd
+ clock_0/gnd clock_0/vdd clock_0/gnd clock_0/vdd clock_0/gnd clock_0/vdd clock_0/gnd
+ clock_0/gnd clock_0/vdd clock_0/gnd clock_0/vdd clock_0/vdd clock_0/vdd clock_0/vdd
+ clock_0/vdd clock_0/vdd clock_0/gnd clock_0/gnd clock_0/gnd clock_0/gnd clock_0/gnd
+ clock_0/vdd clock_0/gnd clock_0/gnd clock_0/vdd clock_0/vdd clock_0/gnd clock_0/vdd
+ clock_0/vdd clock_0/vdd clock_0/vdd clock_0/gnd clock_0/vdd clock_0/gnd clock_0/gnd
+ clock_0/gnd clock_0/gnd clock_0/gnd clock_0/vdd clock_0/vdd clock_0/vdd clock_0/vdd
+ clock_0/gnd clock_0/vdd clock_0/vdd clock_0/vdd clock_0/vdd clock_0/gnd clock_0/vdd
+ clock_0/gnd clock_0/vdd clock_0/vdd clock_0/gnd clock_0/gnd clock_0/vdd clock_0/gnd
+ clock_0/gnd clock_0/vdd clock_0/vdd clock_0/vdd clock_0/gnd clock_0/gnd clock_0/vdd
+ clock_0/gnd clock_0/gnd clock_0/gnd clock_0/vdd clock_0/vdd clock_0/gnd clock_0/vdd
+ clock_0/vdd clock_0/vdd clock_0/gnd clock_0/vdd clock_0/vdd clock_0/gnd clock_0/gnd
+ clock_0/gnd clock_0/vdd clock_0/vdd clock_0/vdd clock_0/gnd clock_0/vdd clock_0/vdd
+ clock_0/vdd clock_0/vdd clock_0/vdd clock_0/vdd clock_0/gnd clock_0/vdd clock_0/gnd
+ clock_0/vdd clock_0/gnd clock_0/gnd clock_0/gnd sky130_fd_pr__nfet_01v8_NJGC8F
Xnmos_diode2_0 out input2 input1 vs nmos_diode2_0/VSUBS nmos_diode2
Xsky130_fd_pr__cap_mim_m3_1_MH6KF8_0 input2 clkb clock_0/gnd sky130_fd_pr__cap_mim_m3_1_MH6KF8
Xsky130_fd_pr__cap_mim_m3_1_MH6KF8_1 input1 clk clock_0/gnd sky130_fd_pr__cap_mim_m3_1_MH6KF8
C0 vs input1 3.39f
C1 clock_0/vdd clkb 17.4f
C2 clock_0/vdd vs 12f
C3 vs clkb 2.33f
C4 input2 input1 8.76f
C5 clock_0/vdd clk 26.5f
C6 vs clk 2.64f
C7 clock_0/vdd out 2.31f
C8 vs out 14.2f
C9 vs input2 4.02f
C10 clock_0/vdd vin 5.36f
C11 vs vin 8.81f
C12 vs nmos_diode2_0/VSUBS 20.1f
C13 out nmos_diode2_0/VSUBS 3.14f
C14 clock_0/a_2432_n962# nmos_diode2_0/VSUBS 8.68f **FLOATING
C15 clock_0/a_2020_n482# nmos_diode2_0/VSUBS 2.57f **FLOATING
C16 clock_0/a_344_102# nmos_diode2_0/VSUBS 2.81f
C17 clock_0/a_2402_572# nmos_diode2_0/VSUBS 2.17f
C18 clock_0/a_344_n986# nmos_diode2_0/VSUBS 2.38f
C19 clock_0/a_3246_118# nmos_diode2_0/VSUBS 6.83f
C20 g2 nmos_diode2_0/VSUBS 2.44f
C21 capacitors_5_0/capacitor_5_4/buffer_and_gate_0/and_gate_0/a_n78_396# nmos_diode2_0/VSUBS 2.34f
C22 capacitors_5_0/capacitor_5_4/buffer_and_gate_0/buffer_0/a_1436_1552# nmos_diode2_0/VSUBS 9.98f
C23 capacitors_5_0/capacitor_5_4/buffer_digital_1/in nmos_diode2_0/VSUBS 2.58f
C24 capacitors_5_0/capacitor_5_3/buffer_and_gate_0/and_gate_0/a_n78_396# nmos_diode2_0/VSUBS 2.34f
C25 capacitors_5_0/capacitor_5_3/buffer_and_gate_0/buffer_0/a_1436_1552# nmos_diode2_0/VSUBS 9.98f
C26 capacitors_5_0/capacitor_5_3/buffer_digital_1/in nmos_diode2_0/VSUBS 2.58f
C27 capacitors_5_0/capacitor_5_2/buffer_and_gate_0/and_gate_0/a_n78_396# nmos_diode2_0/VSUBS 2.34f
C28 capacitors_5_0/capacitor_5_2/buffer_and_gate_0/buffer_0/a_1436_1552# nmos_diode2_0/VSUBS 9.98f
C29 capacitors_5_0/capacitor_5_2/buffer_digital_1/in nmos_diode2_0/VSUBS 2.58f
C30 capacitors_5_0/capacitor_5_1/buffer_and_gate_0/and_gate_0/a_n78_396# nmos_diode2_0/VSUBS 2.34f
C31 capacitors_5_0/capacitor_5_1/buffer_and_gate_0/buffer_0/a_1436_1552# nmos_diode2_0/VSUBS 9.98f
C32 capacitors_5_0/capacitor_5_1/buffer_digital_1/in nmos_diode2_0/VSUBS 2.58f
C33 capacitors_5_0/capacitor_5_0/buffer_and_gate_0/and_gate_0/a_n78_396# nmos_diode2_0/VSUBS 2.34f
C34 capacitors_5_0/capacitor_5_0/buffer_and_gate_0/buffer_0/a_1436_1552# nmos_diode2_0/VSUBS 9.98f
C35 capacitors_5_0/capacitor_5_0/buffer_digital_1/in nmos_diode2_0/VSUBS 2.58f
C36 input1 nmos_diode2_0/VSUBS 16.7f
C37 capacitors_5_0/capacitor_5_7/buffer_and_gate_0/and_gate_0/a_n78_396# nmos_diode2_0/VSUBS 2.34f
C38 clk nmos_diode2_0/VSUBS 85f
C39 clock_0/vdd nmos_diode2_0/VSUBS 0.46p
C40 capacitors_5_0/capacitor_5_7/buffer_and_gate_0/buffer_0/a_1436_1552# nmos_diode2_0/VSUBS 9.98f
C41 capacitors_5_0/capacitor_5_7/buffer_digital_1/in nmos_diode2_0/VSUBS 2.58f
C42 capacitors_5_0/capacitor_5_6/buffer_and_gate_0/and_gate_0/a_n78_396# nmos_diode2_0/VSUBS 2.34f
C43 capacitors_5_0/capacitor_5_6/buffer_and_gate_0/buffer_0/a_1436_1552# nmos_diode2_0/VSUBS 9.98f
C44 capacitors_5_0/capacitor_5_6/buffer_digital_1/in nmos_diode2_0/VSUBS 2.58f
C45 capacitors_5_0/capacitor_5_5/buffer_and_gate_0/and_gate_0/a_n78_396# nmos_diode2_0/VSUBS 2.34f
C46 capacitors_5_0/capacitor_5_5/buffer_and_gate_0/buffer_0/a_1436_1552# nmos_diode2_0/VSUBS 9.98f
C47 capacitors_5_0/capacitor_5_5/buffer_digital_1/in nmos_diode2_0/VSUBS 2.58f
C48 capacitors_5_1/capacitor_5_4/buffer_and_gate_0/and_gate_0/a_n78_396# nmos_diode2_0/VSUBS 2.34f
C49 capacitors_5_1/capacitor_5_4/buffer_and_gate_0/buffer_0/a_1436_1552# nmos_diode2_0/VSUBS 9.98f
C50 capacitors_5_1/capacitor_5_4/buffer_digital_1/in nmos_diode2_0/VSUBS 2.58f
C51 capacitors_5_1/capacitor_5_3/buffer_and_gate_0/and_gate_0/a_n78_396# nmos_diode2_0/VSUBS 2.34f
C52 capacitors_5_1/capacitor_5_3/buffer_and_gate_0/buffer_0/a_1436_1552# nmos_diode2_0/VSUBS 9.98f
C53 capacitors_5_1/capacitor_5_3/buffer_digital_1/in nmos_diode2_0/VSUBS 2.58f
C54 capacitors_5_1/capacitor_5_2/buffer_and_gate_0/and_gate_0/a_n78_396# nmos_diode2_0/VSUBS 2.34f
C55 capacitors_5_1/capacitor_5_2/buffer_and_gate_0/buffer_0/a_1436_1552# nmos_diode2_0/VSUBS 9.98f
C56 capacitors_5_1/capacitor_5_2/buffer_digital_1/in nmos_diode2_0/VSUBS 2.58f
C57 capacitors_5_1/capacitor_5_1/buffer_and_gate_0/and_gate_0/a_n78_396# nmos_diode2_0/VSUBS 2.34f
C58 capacitors_5_1/capacitor_5_1/buffer_and_gate_0/buffer_0/a_1436_1552# nmos_diode2_0/VSUBS 9.98f
C59 capacitors_5_1/capacitor_5_1/buffer_digital_1/in nmos_diode2_0/VSUBS 2.58f
C60 capacitors_5_1/capacitor_5_0/buffer_and_gate_0/and_gate_0/a_n78_396# nmos_diode2_0/VSUBS 2.34f
C61 capacitors_5_1/capacitor_5_0/buffer_and_gate_0/buffer_0/a_1436_1552# nmos_diode2_0/VSUBS 9.98f
C62 capacitors_5_1/capacitor_5_0/buffer_digital_1/in nmos_diode2_0/VSUBS 2.58f
C63 input2 nmos_diode2_0/VSUBS 16.9f
C64 capacitors_5_1/capacitor_5_7/buffer_and_gate_0/and_gate_0/a_n78_396# nmos_diode2_0/VSUBS 2.34f
C65 clkb nmos_diode2_0/VSUBS 87.1f
C66 capacitors_5_1/capacitor_5_7/buffer_and_gate_0/buffer_0/a_1436_1552# nmos_diode2_0/VSUBS 9.98f
C67 capacitors_5_1/capacitor_5_7/buffer_digital_1/in nmos_diode2_0/VSUBS 2.58f
C68 capacitors_5_1/capacitor_5_6/buffer_and_gate_0/and_gate_0/a_n78_396# nmos_diode2_0/VSUBS 2.34f
C69 capacitors_5_1/capacitor_5_6/buffer_and_gate_0/buffer_0/a_1436_1552# nmos_diode2_0/VSUBS 9.98f
C70 capacitors_5_1/capacitor_5_6/buffer_digital_1/in nmos_diode2_0/VSUBS 2.58f
C71 capacitors_5_1/capacitor_5_5/buffer_and_gate_0/and_gate_0/a_n78_396# nmos_diode2_0/VSUBS 2.34f
C72 capacitors_5_1/capacitor_5_5/buffer_and_gate_0/buffer_0/a_1436_1552# nmos_diode2_0/VSUBS 9.98f
C73 capacitors_5_1/capacitor_5_5/buffer_digital_1/in nmos_diode2_0/VSUBS 2.58f
C74 g1 nmos_diode2_0/VSUBS 2.64f
.ends

.subckt cp2_buffer1 charge_pump_0/a_18057_18271# charge_pump_0/in4 buffer_digital_0/in
+ charge_pump_0/in5 charge_pump_0/vin charge_pump_0/out charge_pump_0/in6 charge_pump_0/in7
+ charge_pump_0/vs charge_pump_0/in8 charge_pump_0/in1 charge_pump_0/in3 charge_pump_0/in2
+ buffer_digital_1/i VSUBS buffer_digital_1/VDD
Xpmos_decap_10_10 VSUBS buffer_digital_1/VDD VSUBS pmos_decap_10
Xpmos_decap_10_11 VSUBS buffer_digital_1/VDD VSUBS pmos_decap_10
Xpmos_decap_10_12 VSUBS buffer_digital_1/VDD VSUBS pmos_decap_10
Xpmos_decap_10_13 VSUBS buffer_digital_1/VDD VSUBS pmos_decap_10
Xcharge_pump_0 charge_pump_0/in1 charge_pump_0/in3 charge_pump_0/in5 charge_pump_0/input1
+ charge_pump_0/input2 charge_pump_0/out charge_pump_0/clk charge_pump_0/clkb buffer_digital_0/in
+ charge_pump_0/g1 charge_pump_0/g2 charge_pump_0/vin charge_pump_0/a_18057_18271#
+ charge_pump_0/in6 charge_pump_0/in8 charge_pump_0/in4 charge_pump_0/in7 charge_pump_0/in2
+ charge_pump_0/vs VSUBS buffer_digital_1/VDD charge_pump
Xbuffer_digital_0 buffer_digital_0/i buffer_digital_0/in buffer_digital_1/VDD VSUBS
+ buffer_digital
Xbuffer_digital_1 buffer_digital_1/i buffer_digital_0/i buffer_digital_1/VDD VSUBS
+ buffer_digital
Xnmos_decap_10_0 buffer_digital_1/VDD VSUBS VSUBS nmos_decap_10
Xnmos_decap_10_1 buffer_digital_1/VDD VSUBS VSUBS nmos_decap_10
Xnmos_decap_10_2 buffer_digital_1/VDD VSUBS VSUBS nmos_decap_10
Xnmos_decap_10_3 buffer_digital_1/VDD VSUBS VSUBS nmos_decap_10
Xnmos_decap_10_4 buffer_digital_1/VDD VSUBS VSUBS nmos_decap_10
Xnmos_decap_10_5 buffer_digital_1/VDD VSUBS VSUBS nmos_decap_10
Xpmos_decap_10_0 VSUBS buffer_digital_1/VDD VSUBS pmos_decap_10
Xpmos_decap_10_1 VSUBS buffer_digital_1/VDD VSUBS pmos_decap_10
Xpmos_decap_10_2 VSUBS buffer_digital_1/VDD VSUBS pmos_decap_10
Xpmos_decap_10_3 VSUBS buffer_digital_1/VDD VSUBS pmos_decap_10
Xpmos_decap_10_4 VSUBS buffer_digital_1/VDD VSUBS pmos_decap_10
Xpmos_decap_10_5 VSUBS buffer_digital_1/VDD VSUBS pmos_decap_10
Xpmos_decap_10_6 VSUBS buffer_digital_1/VDD VSUBS pmos_decap_10
Xpmos_decap_10_7 VSUBS buffer_digital_1/VDD VSUBS pmos_decap_10
Xpmos_decap_10_9 VSUBS buffer_digital_1/VDD VSUBS pmos_decap_10
Xpmos_decap_10_8 VSUBS buffer_digital_1/VDD VSUBS pmos_decap_10
C0 buffer_digital_1/VDD buffer_digital_0/in 4.8f
C1 buffer_digital_1/VDD buffer_digital_1/i 3.74f
C2 buffer_digital_1/i charge_pump_0/nmos_diode2_0/VSUBS 8.29f
C3 charge_pump_0/vs charge_pump_0/nmos_diode2_0/VSUBS 19f
C4 charge_pump_0/clock_0/a_2432_n962# charge_pump_0/nmos_diode2_0/VSUBS 8.68f **FLOATING
C5 charge_pump_0/clock_0/a_2020_n482# charge_pump_0/nmos_diode2_0/VSUBS 2.57f **FLOATING
C6 charge_pump_0/clock_0/a_344_102# charge_pump_0/nmos_diode2_0/VSUBS 2.81f
C7 charge_pump_0/clock_0/a_2402_572# charge_pump_0/nmos_diode2_0/VSUBS 2.17f
C8 charge_pump_0/clock_0/a_344_n986# charge_pump_0/nmos_diode2_0/VSUBS 2.38f
C9 buffer_digital_0/in charge_pump_0/nmos_diode2_0/VSUBS 12.9f
C10 charge_pump_0/clock_0/a_3246_118# charge_pump_0/nmos_diode2_0/VSUBS 6.83f
C11 charge_pump_0/g2 charge_pump_0/nmos_diode2_0/VSUBS 2.44f
C12 charge_pump_0/capacitors_5_0/capacitor_5_4/buffer_and_gate_0/and_gate_0/a_n78_396# charge_pump_0/nmos_diode2_0/VSUBS 2.34f
C13 charge_pump_0/capacitors_5_0/capacitor_5_4/buffer_and_gate_0/buffer_0/a_1436_1552# charge_pump_0/nmos_diode2_0/VSUBS 9.98f
C14 charge_pump_0/capacitors_5_0/capacitor_5_4/buffer_digital_1/in charge_pump_0/nmos_diode2_0/VSUBS 2.58f
C15 charge_pump_0/capacitors_5_0/capacitor_5_3/buffer_and_gate_0/and_gate_0/a_n78_396# charge_pump_0/nmos_diode2_0/VSUBS 2.34f
C16 charge_pump_0/capacitors_5_0/capacitor_5_3/buffer_and_gate_0/buffer_0/a_1436_1552# charge_pump_0/nmos_diode2_0/VSUBS 9.98f
C17 charge_pump_0/capacitors_5_0/capacitor_5_3/buffer_digital_1/in charge_pump_0/nmos_diode2_0/VSUBS 2.58f
C18 charge_pump_0/capacitors_5_0/capacitor_5_2/buffer_and_gate_0/and_gate_0/a_n78_396# charge_pump_0/nmos_diode2_0/VSUBS 2.34f
C19 charge_pump_0/capacitors_5_0/capacitor_5_2/buffer_and_gate_0/buffer_0/a_1436_1552# charge_pump_0/nmos_diode2_0/VSUBS 9.98f
C20 charge_pump_0/capacitors_5_0/capacitor_5_2/buffer_digital_1/in charge_pump_0/nmos_diode2_0/VSUBS 2.58f
C21 charge_pump_0/capacitors_5_0/capacitor_5_1/buffer_and_gate_0/and_gate_0/a_n78_396# charge_pump_0/nmos_diode2_0/VSUBS 2.34f
C22 charge_pump_0/capacitors_5_0/capacitor_5_1/buffer_and_gate_0/buffer_0/a_1436_1552# charge_pump_0/nmos_diode2_0/VSUBS 9.98f
C23 charge_pump_0/capacitors_5_0/capacitor_5_1/buffer_digital_1/in charge_pump_0/nmos_diode2_0/VSUBS 2.58f
C24 charge_pump_0/capacitors_5_0/capacitor_5_0/buffer_and_gate_0/and_gate_0/a_n78_396# charge_pump_0/nmos_diode2_0/VSUBS 2.34f
C25 charge_pump_0/capacitors_5_0/capacitor_5_0/buffer_and_gate_0/buffer_0/a_1436_1552# charge_pump_0/nmos_diode2_0/VSUBS 9.98f
C26 charge_pump_0/capacitors_5_0/capacitor_5_0/buffer_digital_1/in charge_pump_0/nmos_diode2_0/VSUBS 2.58f
C27 charge_pump_0/input1 charge_pump_0/nmos_diode2_0/VSUBS 15f
C28 charge_pump_0/capacitors_5_0/capacitor_5_7/buffer_and_gate_0/and_gate_0/a_n78_396# charge_pump_0/nmos_diode2_0/VSUBS 2.34f
C29 charge_pump_0/clk charge_pump_0/nmos_diode2_0/VSUBS 82.8f
C30 buffer_digital_1/VDD charge_pump_0/nmos_diode2_0/VSUBS 0.525p
C31 charge_pump_0/capacitors_5_0/capacitor_5_7/buffer_and_gate_0/buffer_0/a_1436_1552# charge_pump_0/nmos_diode2_0/VSUBS 9.98f
C32 charge_pump_0/capacitors_5_0/capacitor_5_7/buffer_digital_1/in charge_pump_0/nmos_diode2_0/VSUBS 2.58f
C33 charge_pump_0/capacitors_5_0/capacitor_5_6/buffer_and_gate_0/and_gate_0/a_n78_396# charge_pump_0/nmos_diode2_0/VSUBS 2.34f
C34 charge_pump_0/capacitors_5_0/capacitor_5_6/buffer_and_gate_0/buffer_0/a_1436_1552# charge_pump_0/nmos_diode2_0/VSUBS 9.98f
C35 charge_pump_0/capacitors_5_0/capacitor_5_6/buffer_digital_1/in charge_pump_0/nmos_diode2_0/VSUBS 2.58f
C36 charge_pump_0/capacitors_5_0/capacitor_5_5/buffer_and_gate_0/and_gate_0/a_n78_396# charge_pump_0/nmos_diode2_0/VSUBS 2.34f
C37 charge_pump_0/capacitors_5_0/capacitor_5_5/buffer_and_gate_0/buffer_0/a_1436_1552# charge_pump_0/nmos_diode2_0/VSUBS 9.98f
C38 charge_pump_0/capacitors_5_0/capacitor_5_5/buffer_digital_1/in charge_pump_0/nmos_diode2_0/VSUBS 2.58f
C39 charge_pump_0/capacitors_5_1/capacitor_5_4/buffer_and_gate_0/and_gate_0/a_n78_396# charge_pump_0/nmos_diode2_0/VSUBS 2.34f
C40 charge_pump_0/capacitors_5_1/capacitor_5_4/buffer_and_gate_0/buffer_0/a_1436_1552# charge_pump_0/nmos_diode2_0/VSUBS 9.98f
C41 charge_pump_0/capacitors_5_1/capacitor_5_4/buffer_digital_1/in charge_pump_0/nmos_diode2_0/VSUBS 2.58f
C42 charge_pump_0/capacitors_5_1/capacitor_5_3/buffer_and_gate_0/and_gate_0/a_n78_396# charge_pump_0/nmos_diode2_0/VSUBS 2.34f
C43 charge_pump_0/capacitors_5_1/capacitor_5_3/buffer_and_gate_0/buffer_0/a_1436_1552# charge_pump_0/nmos_diode2_0/VSUBS 9.98f
C44 charge_pump_0/capacitors_5_1/capacitor_5_3/buffer_digital_1/in charge_pump_0/nmos_diode2_0/VSUBS 2.58f
C45 charge_pump_0/capacitors_5_1/capacitor_5_2/buffer_and_gate_0/and_gate_0/a_n78_396# charge_pump_0/nmos_diode2_0/VSUBS 2.34f
C46 charge_pump_0/capacitors_5_1/capacitor_5_2/buffer_and_gate_0/buffer_0/a_1436_1552# charge_pump_0/nmos_diode2_0/VSUBS 9.98f
C47 charge_pump_0/capacitors_5_1/capacitor_5_2/buffer_digital_1/in charge_pump_0/nmos_diode2_0/VSUBS 2.58f
C48 charge_pump_0/capacitors_5_1/capacitor_5_1/buffer_and_gate_0/and_gate_0/a_n78_396# charge_pump_0/nmos_diode2_0/VSUBS 2.34f
C49 charge_pump_0/capacitors_5_1/capacitor_5_1/buffer_and_gate_0/buffer_0/a_1436_1552# charge_pump_0/nmos_diode2_0/VSUBS 9.98f
C50 charge_pump_0/capacitors_5_1/capacitor_5_1/buffer_digital_1/in charge_pump_0/nmos_diode2_0/VSUBS 2.58f
C51 charge_pump_0/capacitors_5_1/capacitor_5_0/buffer_and_gate_0/and_gate_0/a_n78_396# charge_pump_0/nmos_diode2_0/VSUBS 2.34f
C52 charge_pump_0/capacitors_5_1/capacitor_5_0/buffer_and_gate_0/buffer_0/a_1436_1552# charge_pump_0/nmos_diode2_0/VSUBS 9.98f
C53 charge_pump_0/capacitors_5_1/capacitor_5_0/buffer_digital_1/in charge_pump_0/nmos_diode2_0/VSUBS 2.58f
C54 charge_pump_0/input2 charge_pump_0/nmos_diode2_0/VSUBS 14.4f
C55 charge_pump_0/capacitors_5_1/capacitor_5_7/buffer_and_gate_0/and_gate_0/a_n78_396# charge_pump_0/nmos_diode2_0/VSUBS 2.34f
C56 charge_pump_0/clkb charge_pump_0/nmos_diode2_0/VSUBS 83.9f
C57 charge_pump_0/capacitors_5_1/capacitor_5_7/buffer_and_gate_0/buffer_0/a_1436_1552# charge_pump_0/nmos_diode2_0/VSUBS 9.98f
C58 charge_pump_0/capacitors_5_1/capacitor_5_7/buffer_digital_1/in charge_pump_0/nmos_diode2_0/VSUBS 2.58f
C59 charge_pump_0/capacitors_5_1/capacitor_5_6/buffer_and_gate_0/and_gate_0/a_n78_396# charge_pump_0/nmos_diode2_0/VSUBS 2.34f
C60 charge_pump_0/capacitors_5_1/capacitor_5_6/buffer_and_gate_0/buffer_0/a_1436_1552# charge_pump_0/nmos_diode2_0/VSUBS 9.98f
C61 charge_pump_0/capacitors_5_1/capacitor_5_6/buffer_digital_1/in charge_pump_0/nmos_diode2_0/VSUBS 2.58f
C62 charge_pump_0/capacitors_5_1/capacitor_5_5/buffer_and_gate_0/and_gate_0/a_n78_396# charge_pump_0/nmos_diode2_0/VSUBS 2.34f
C63 charge_pump_0/capacitors_5_1/capacitor_5_5/buffer_and_gate_0/buffer_0/a_1436_1552# charge_pump_0/nmos_diode2_0/VSUBS 9.98f
C64 charge_pump_0/capacitors_5_1/capacitor_5_5/buffer_digital_1/in charge_pump_0/nmos_diode2_0/VSUBS 2.58f
C65 charge_pump_0/g1 charge_pump_0/nmos_diode2_0/VSUBS 2.63f
.ends

.subckt charge_pump_reverse m1_11946_n452# nmos_dnw3_0/vin capacitors_5_1/capacitor_5_2/i1
+ capacitors_5_1/capacitor_5_3/i1 a_18057_18271# capacitors_5_1/capacitor_5_4/i1 capacitors_5_1/capacitor_5_5/i1
+ clock_0/clk_in clock_0/vdd capacitors_5_1/capacitor_5_0/i1 capacitors_5_1/capacitor_5_7/i1
+ clock_0/gnd capacitors_5_1/capacitor_5_6/i1 capacitors_5_1/capacitor_5_1/i1 nmos_dnw3_0/vs
Xsky130_fd_pr__cap_mim_m3_1_MH6KF8_4 nmos_dnw3_0/clk clock_0/clkb clock_0/gnd sky130_fd_pr__cap_mim_m3_1_MH6KF8
Xsky130_fd_pr__cap_mim_m3_1_MH6KF8_5 nmos_dnw3_0/clkb clock_0/clk clock_0/gnd sky130_fd_pr__cap_mim_m3_1_MH6KF8
Xcapacitors_5_1 capacitors_5_1/capacitor_5_7/i1 capacitors_5_1/capacitor_5_1/i1 capacitors_5_1/capacitor_5_6/i1
+ capacitors_5_1/capacitor_5_0/i1 clock_0/vdd capacitors_5_1/capacitor_5_3/i1 clock_0/vdd
+ clock_0/vdd nmos_dnw3_0/out2 capacitors_5_1/capacitor_5_4/i1 capacitors_5_1/capacitor_5_2/i1
+ clock_0/clk clock_0/vdd capacitors_5_1/capacitor_5_5/i1 clock_0/gnd clock_0/vdd
+ capacitors_5
Xcapacitors_5_0 capacitors_5_1/capacitor_5_7/i1 capacitors_5_1/capacitor_5_1/i1 capacitors_5_1/capacitor_5_6/i1
+ capacitors_5_1/capacitor_5_0/i1 clock_0/vdd capacitors_5_1/capacitor_5_3/i1 clock_0/vdd
+ clock_0/vdd nmos_dnw3_0/out1 capacitors_5_1/capacitor_5_4/i1 capacitors_5_1/capacitor_5_2/i1
+ clock_0/clkb clock_0/vdd capacitors_5_1/capacitor_5_5/i1 clock_0/gnd clock_0/vdd
+ capacitors_5
Xnmos_dnw3_0 nmos_dnw3_0/vin nmos_dnw3_0/out1 nmos_dnw3_0/out2 nmos_dnw3_0/clk nmos_dnw3_0/clkb
+ nmos_dnw3_0/vs clock_0/gnd nmos_dnw3
Xclock_0 clock_0/clk_in clock_0/vdd clock_0/gnd clock_0/clk clock_0/clkb clock
Xsky130_fd_pr__pfet_01v8_4RPJ49_0 clock_0/gnd clock_0/vdd clock_0/vdd clock_0/gnd
+ clock_0/gnd clock_0/vdd clock_0/vdd clock_0/vdd clock_0/gnd clock_0/vdd clock_0/gnd
+ clock_0/gnd clock_0/vdd clock_0/gnd clock_0/gnd clock_0/gnd clock_0/vdd clock_0/vdd
+ clock_0/vdd clock_0/vdd clock_0/gnd clock_0/vdd clock_0/gnd clock_0/gnd clock_0/gnd
+ clock_0/gnd clock_0/gnd clock_0/gnd clock_0/gnd clock_0/vdd clock_0/gnd clock_0/vdd
+ clock_0/gnd clock_0/gnd clock_0/vdd clock_0/gnd clock_0/gnd clock_0/vdd clock_0/vdd
+ clock_0/gnd clock_0/vdd clock_0/gnd clock_0/gnd clock_0/vdd clock_0/gnd clock_0/gnd
+ clock_0/vdd clock_0/vdd clock_0/gnd clock_0/gnd clock_0/vdd clock_0/vdd clock_0/vdd
+ clock_0/gnd clock_0/gnd clock_0/vdd clock_0/vdd clock_0/gnd clock_0/gnd clock_0/vdd
+ clock_0/vdd clock_0/gnd clock_0/vdd clock_0/gnd clock_0/vdd clock_0/gnd clock_0/gnd
+ clock_0/gnd clock_0/vdd clock_0/gnd clock_0/gnd clock_0/gnd clock_0/vdd clock_0/vdd
+ clock_0/gnd clock_0/gnd clock_0/vdd clock_0/vdd clock_0/gnd clock_0/gnd clock_0/vdd
+ clock_0/vdd clock_0/gnd clock_0/gnd clock_0/gnd clock_0/vdd clock_0/vdd clock_0/vdd
+ clock_0/vdd clock_0/vdd clock_0/vdd clock_0/vdd clock_0/vdd clock_0/vdd clock_0/gnd
+ clock_0/gnd clock_0/vdd clock_0/vdd clock_0/vdd clock_0/gnd clock_0/vdd clock_0/vdd
+ clock_0/vdd clock_0/vdd clock_0/vdd clock_0/gnd clock_0/vdd clock_0/vdd clock_0/gnd
+ clock_0/vdd clock_0/vdd clock_0/gnd clock_0/gnd clock_0/gnd clock_0/gnd clock_0/gnd
+ clock_0/vdd clock_0/vdd clock_0/vdd clock_0/gnd clock_0/vdd clock_0/vdd clock_0/gnd
+ clock_0/vdd clock_0/gnd clock_0/vdd clock_0/vdd clock_0/vdd clock_0/gnd clock_0/gnd
+ clock_0/vdd clock_0/vdd clock_0/gnd clock_0/vdd clock_0/vdd clock_0/vdd clock_0/vdd
+ clock_0/gnd clock_0/vdd clock_0/gnd clock_0/gnd clock_0/gnd clock_0/vdd clock_0/vdd
+ clock_0/vdd clock_0/gnd clock_0/gnd clock_0/gnd clock_0/gnd clock_0/vdd clock_0/gnd
+ clock_0/gnd clock_0/gnd clock_0/vdd clock_0/gnd clock_0/gnd clock_0/gnd clock_0/gnd
+ clock_0/vdd clock_0/gnd clock_0/gnd clock_0/vdd clock_0/vdd sky130_fd_pr__pfet_01v8_4RPJ49
Xsky130_fd_pr__pfet_01v8_4RPJ49_1 clock_0/gnd clock_0/vdd clock_0/vdd clock_0/gnd
+ clock_0/gnd clock_0/vdd clock_0/vdd clock_0/vdd clock_0/gnd clock_0/vdd clock_0/gnd
+ clock_0/gnd clock_0/vdd clock_0/gnd clock_0/gnd clock_0/gnd clock_0/vdd clock_0/vdd
+ clock_0/vdd clock_0/vdd clock_0/gnd clock_0/vdd clock_0/gnd clock_0/gnd clock_0/gnd
+ clock_0/gnd clock_0/gnd clock_0/gnd clock_0/gnd clock_0/vdd clock_0/gnd clock_0/vdd
+ clock_0/gnd clock_0/gnd clock_0/vdd clock_0/gnd clock_0/gnd clock_0/vdd clock_0/vdd
+ clock_0/gnd clock_0/vdd clock_0/gnd clock_0/gnd clock_0/vdd clock_0/gnd clock_0/gnd
+ clock_0/vdd clock_0/vdd clock_0/gnd clock_0/gnd clock_0/vdd clock_0/vdd clock_0/vdd
+ clock_0/gnd clock_0/gnd clock_0/vdd clock_0/vdd clock_0/gnd clock_0/gnd clock_0/vdd
+ clock_0/vdd clock_0/gnd clock_0/vdd clock_0/gnd clock_0/vdd clock_0/gnd clock_0/gnd
+ clock_0/gnd clock_0/vdd clock_0/gnd clock_0/gnd clock_0/gnd clock_0/vdd clock_0/vdd
+ clock_0/gnd clock_0/gnd clock_0/vdd clock_0/vdd clock_0/gnd clock_0/gnd clock_0/vdd
+ clock_0/vdd clock_0/gnd clock_0/gnd clock_0/gnd clock_0/vdd clock_0/vdd clock_0/vdd
+ clock_0/vdd clock_0/vdd clock_0/vdd clock_0/vdd clock_0/vdd clock_0/vdd clock_0/gnd
+ clock_0/gnd clock_0/vdd clock_0/vdd clock_0/vdd clock_0/gnd clock_0/vdd clock_0/vdd
+ clock_0/vdd clock_0/vdd clock_0/vdd clock_0/gnd clock_0/vdd clock_0/vdd clock_0/gnd
+ clock_0/vdd clock_0/vdd clock_0/gnd clock_0/gnd clock_0/gnd clock_0/gnd clock_0/gnd
+ clock_0/vdd clock_0/vdd clock_0/vdd clock_0/gnd clock_0/vdd clock_0/vdd clock_0/gnd
+ clock_0/vdd clock_0/gnd clock_0/vdd clock_0/vdd clock_0/vdd clock_0/gnd clock_0/gnd
+ clock_0/vdd clock_0/vdd clock_0/gnd clock_0/vdd clock_0/vdd clock_0/vdd clock_0/vdd
+ clock_0/gnd clock_0/vdd clock_0/gnd clock_0/gnd clock_0/gnd clock_0/vdd clock_0/vdd
+ clock_0/vdd clock_0/gnd clock_0/gnd clock_0/gnd clock_0/gnd clock_0/vdd clock_0/gnd
+ clock_0/gnd clock_0/gnd clock_0/vdd clock_0/gnd clock_0/gnd clock_0/gnd clock_0/gnd
+ clock_0/vdd clock_0/gnd clock_0/gnd clock_0/vdd clock_0/vdd sky130_fd_pr__pfet_01v8_4RPJ49
Xsky130_fd_pr__nfet_01v8_NJGC8F_0 clock_0/vdd clock_0/gnd clock_0/gnd clock_0/vdd
+ clock_0/vdd clock_0/gnd clock_0/gnd clock_0/vdd clock_0/gnd clock_0/vdd clock_0/gnd
+ clock_0/gnd clock_0/vdd clock_0/gnd clock_0/gnd clock_0/gnd clock_0/vdd clock_0/gnd
+ clock_0/vdd clock_0/vdd clock_0/gnd clock_0/vdd clock_0/vdd clock_0/vdd clock_0/vdd
+ clock_0/gnd clock_0/vdd clock_0/vdd clock_0/gnd clock_0/vdd clock_0/vdd clock_0/gnd
+ clock_0/gnd clock_0/gnd clock_0/gnd clock_0/gnd clock_0/vdd clock_0/gnd clock_0/gnd
+ clock_0/vdd clock_0/gnd clock_0/gnd clock_0/gnd clock_0/vdd clock_0/gnd clock_0/gnd
+ clock_0/vdd clock_0/gnd clock_0/gnd clock_0/gnd clock_0/vdd clock_0/vdd clock_0/gnd
+ clock_0/gnd clock_0/vdd clock_0/gnd clock_0/gnd clock_0/vdd clock_0/gnd clock_0/gnd
+ clock_0/gnd clock_0/vdd clock_0/vdd clock_0/vdd clock_0/gnd clock_0/gnd clock_0/gnd
+ clock_0/gnd clock_0/vdd clock_0/gnd clock_0/vdd clock_0/gnd clock_0/vdd clock_0/gnd
+ clock_0/gnd clock_0/vdd clock_0/gnd clock_0/vdd clock_0/vdd clock_0/vdd clock_0/vdd
+ clock_0/vdd clock_0/vdd clock_0/gnd clock_0/gnd clock_0/gnd clock_0/gnd clock_0/gnd
+ clock_0/vdd clock_0/gnd clock_0/gnd clock_0/vdd clock_0/vdd clock_0/gnd clock_0/vdd
+ clock_0/vdd clock_0/vdd clock_0/vdd clock_0/gnd clock_0/vdd clock_0/gnd clock_0/gnd
+ clock_0/gnd clock_0/gnd clock_0/gnd clock_0/vdd clock_0/vdd clock_0/vdd clock_0/vdd
+ clock_0/gnd clock_0/vdd clock_0/vdd clock_0/vdd clock_0/vdd clock_0/gnd clock_0/vdd
+ clock_0/gnd clock_0/vdd clock_0/vdd clock_0/gnd clock_0/gnd clock_0/vdd clock_0/gnd
+ clock_0/gnd clock_0/vdd clock_0/vdd clock_0/vdd clock_0/gnd clock_0/gnd clock_0/vdd
+ clock_0/gnd clock_0/gnd clock_0/gnd clock_0/vdd clock_0/vdd clock_0/gnd clock_0/vdd
+ clock_0/vdd clock_0/vdd clock_0/gnd clock_0/vdd clock_0/vdd clock_0/gnd clock_0/gnd
+ clock_0/gnd clock_0/vdd clock_0/vdd clock_0/vdd clock_0/gnd clock_0/vdd clock_0/vdd
+ clock_0/vdd clock_0/vdd clock_0/vdd clock_0/vdd clock_0/gnd clock_0/vdd clock_0/gnd
+ clock_0/vdd clock_0/gnd clock_0/gnd clock_0/gnd sky130_fd_pr__nfet_01v8_NJGC8F
Xsky130_fd_pr__nfet_01v8_NJGC8F_1 clock_0/vdd clock_0/gnd clock_0/gnd clock_0/vdd
+ clock_0/vdd clock_0/gnd clock_0/gnd clock_0/vdd clock_0/gnd clock_0/vdd clock_0/gnd
+ clock_0/gnd clock_0/vdd clock_0/gnd clock_0/gnd clock_0/gnd clock_0/vdd clock_0/gnd
+ clock_0/vdd clock_0/vdd clock_0/gnd clock_0/vdd clock_0/vdd clock_0/vdd clock_0/vdd
+ clock_0/gnd clock_0/vdd clock_0/vdd clock_0/gnd clock_0/vdd clock_0/vdd clock_0/gnd
+ clock_0/gnd clock_0/gnd clock_0/gnd clock_0/gnd clock_0/vdd clock_0/gnd clock_0/gnd
+ clock_0/vdd clock_0/gnd clock_0/gnd clock_0/gnd clock_0/vdd clock_0/gnd clock_0/gnd
+ clock_0/vdd clock_0/gnd clock_0/gnd clock_0/gnd clock_0/vdd clock_0/vdd clock_0/gnd
+ clock_0/gnd clock_0/vdd clock_0/gnd clock_0/gnd clock_0/vdd clock_0/gnd clock_0/gnd
+ clock_0/gnd clock_0/vdd clock_0/vdd clock_0/vdd clock_0/gnd clock_0/gnd clock_0/gnd
+ clock_0/gnd clock_0/vdd clock_0/gnd clock_0/vdd clock_0/gnd clock_0/vdd clock_0/gnd
+ clock_0/gnd clock_0/vdd clock_0/gnd clock_0/vdd clock_0/vdd clock_0/vdd clock_0/vdd
+ clock_0/vdd clock_0/vdd clock_0/gnd clock_0/gnd clock_0/gnd clock_0/gnd clock_0/gnd
+ clock_0/vdd clock_0/gnd clock_0/gnd clock_0/vdd clock_0/vdd clock_0/gnd clock_0/vdd
+ clock_0/vdd clock_0/vdd clock_0/vdd clock_0/gnd clock_0/vdd clock_0/gnd clock_0/gnd
+ clock_0/gnd clock_0/gnd clock_0/gnd clock_0/vdd clock_0/vdd clock_0/vdd clock_0/vdd
+ clock_0/gnd clock_0/vdd clock_0/vdd clock_0/vdd clock_0/vdd clock_0/gnd clock_0/vdd
+ clock_0/gnd clock_0/vdd clock_0/vdd clock_0/gnd clock_0/gnd clock_0/vdd clock_0/gnd
+ clock_0/gnd clock_0/vdd clock_0/vdd clock_0/vdd clock_0/gnd clock_0/gnd clock_0/vdd
+ clock_0/gnd clock_0/gnd clock_0/gnd clock_0/vdd clock_0/vdd clock_0/gnd clock_0/vdd
+ clock_0/vdd clock_0/vdd clock_0/gnd clock_0/vdd clock_0/vdd clock_0/gnd clock_0/gnd
+ clock_0/gnd clock_0/vdd clock_0/vdd clock_0/vdd clock_0/gnd clock_0/vdd clock_0/vdd
+ clock_0/vdd clock_0/vdd clock_0/vdd clock_0/vdd clock_0/gnd clock_0/vdd clock_0/gnd
+ clock_0/vdd clock_0/gnd clock_0/gnd clock_0/gnd sky130_fd_pr__nfet_01v8_NJGC8F
Xnmos_diode2_0 m1_11946_n452# nmos_dnw3_0/out2 nmos_dnw3_0/out1 nmos_dnw3_0/vs clock_0/gnd
+ nmos_diode2
Xsky130_fd_pr__cap_mim_m3_1_MH6KF8_0 nmos_dnw3_0/out2 clock_0/clk clock_0/gnd sky130_fd_pr__cap_mim_m3_1_MH6KF8
Xsky130_fd_pr__cap_mim_m3_1_MH6KF8_1 nmos_dnw3_0/out1 clock_0/clkb clock_0/gnd sky130_fd_pr__cap_mim_m3_1_MH6KF8
C0 nmos_dnw3_0/out1 nmos_dnw3_0/out2 8.76f
C1 nmos_dnw3_0/out1 nmos_dnw3_0/vs 3.31f
C2 nmos_dnw3_0/out2 nmos_dnw3_0/vs 5.26f
C3 clock_0/vdd nmos_dnw3_0/vs 2.47f
C4 clock_0/clk clock_0/vdd 20f
C5 clock_0/vdd nmos_dnw3_0/vin 8.88f
C6 m1_11946_n452# nmos_dnw3_0/vs 13.5f
C7 m1_11946_n452# clock_0/vdd 2.54f
C8 clock_0/vdd clock_0/clkb 24.4f
C9 nmos_dnw3_0/vs clock_0/gnd 19.5f
C10 m1_11946_n452# clock_0/gnd 2.97f
C11 clock_0/a_2432_n962# clock_0/gnd 8.69f **FLOATING
C12 clock_0/a_2020_n482# clock_0/gnd 2.57f **FLOATING
C13 clock_0/a_344_102# clock_0/gnd 2.81f
C14 clock_0/a_2402_572# clock_0/gnd 2.17f
C15 clock_0/a_344_n986# clock_0/gnd 2.38f
C16 clock_0/a_3246_118# clock_0/gnd 6.83f
C17 nmos_dnw3_0/vin clock_0/gnd 2.5f
C18 nmos_dnw3_0/clkb clock_0/gnd 2.24f
C19 capacitors_5_0/capacitor_5_4/buffer_and_gate_0/and_gate_0/a_n78_396# clock_0/gnd 2.34f
C20 capacitors_5_0/capacitor_5_4/buffer_and_gate_0/buffer_0/a_1436_1552# clock_0/gnd 9.98f
C21 capacitors_5_0/capacitor_5_4/buffer_digital_1/in clock_0/gnd 2.58f
C22 capacitors_5_0/capacitor_5_3/buffer_and_gate_0/and_gate_0/a_n78_396# clock_0/gnd 2.34f
C23 capacitors_5_0/capacitor_5_3/buffer_and_gate_0/buffer_0/a_1436_1552# clock_0/gnd 9.98f
C24 capacitors_5_0/capacitor_5_3/buffer_digital_1/in clock_0/gnd 2.58f
C25 capacitors_5_0/capacitor_5_2/buffer_and_gate_0/and_gate_0/a_n78_396# clock_0/gnd 2.34f
C26 capacitors_5_0/capacitor_5_2/buffer_and_gate_0/buffer_0/a_1436_1552# clock_0/gnd 9.98f
C27 capacitors_5_0/capacitor_5_2/buffer_digital_1/in clock_0/gnd 2.58f
C28 capacitors_5_0/capacitor_5_1/buffer_and_gate_0/and_gate_0/a_n78_396# clock_0/gnd 2.34f
C29 capacitors_5_0/capacitor_5_1/buffer_and_gate_0/buffer_0/a_1436_1552# clock_0/gnd 9.98f
C30 capacitors_5_0/capacitor_5_1/buffer_digital_1/in clock_0/gnd 2.58f
C31 capacitors_5_0/capacitor_5_0/buffer_and_gate_0/and_gate_0/a_n78_396# clock_0/gnd 2.34f
C32 capacitors_5_0/capacitor_5_0/buffer_and_gate_0/buffer_0/a_1436_1552# clock_0/gnd 9.98f
C33 capacitors_5_0/capacitor_5_0/buffer_digital_1/in clock_0/gnd 2.58f
C34 nmos_dnw3_0/out1 clock_0/gnd 16.7f
C35 capacitors_5_0/capacitor_5_7/buffer_and_gate_0/and_gate_0/a_n78_396# clock_0/gnd 2.34f
C36 clock_0/clkb clock_0/gnd 92.4f
C37 capacitors_5_0/capacitor_5_7/buffer_and_gate_0/buffer_0/a_1436_1552# clock_0/gnd 9.98f
C38 capacitors_5_0/capacitor_5_7/buffer_digital_1/in clock_0/gnd 2.58f
C39 capacitors_5_0/capacitor_5_6/buffer_and_gate_0/and_gate_0/a_n78_396# clock_0/gnd 2.34f
C40 capacitors_5_0/capacitor_5_6/buffer_and_gate_0/buffer_0/a_1436_1552# clock_0/gnd 9.98f
C41 capacitors_5_0/capacitor_5_6/buffer_digital_1/in clock_0/gnd 2.58f
C42 capacitors_5_0/capacitor_5_5/buffer_and_gate_0/and_gate_0/a_n78_396# clock_0/gnd 2.34f
C43 capacitors_5_0/capacitor_5_5/buffer_and_gate_0/buffer_0/a_1436_1552# clock_0/gnd 9.98f
C44 capacitors_5_0/capacitor_5_5/buffer_digital_1/in clock_0/gnd 2.58f
C45 capacitors_5_1/capacitor_5_4/buffer_and_gate_0/and_gate_0/a_n78_396# clock_0/gnd 2.34f
C46 capacitors_5_1/capacitor_5_4/buffer_and_gate_0/buffer_0/a_1436_1552# clock_0/gnd 9.98f
C47 capacitors_5_1/capacitor_5_4/buffer_digital_1/in clock_0/gnd 2.58f
C48 capacitors_5_1/capacitor_5_3/buffer_and_gate_0/and_gate_0/a_n78_396# clock_0/gnd 2.34f
C49 capacitors_5_1/capacitor_5_3/buffer_and_gate_0/buffer_0/a_1436_1552# clock_0/gnd 9.98f
C50 capacitors_5_1/capacitor_5_3/buffer_digital_1/in clock_0/gnd 2.58f
C51 capacitors_5_1/capacitor_5_2/buffer_and_gate_0/and_gate_0/a_n78_396# clock_0/gnd 2.34f
C52 capacitors_5_1/capacitor_5_2/buffer_and_gate_0/buffer_0/a_1436_1552# clock_0/gnd 9.98f
C53 capacitors_5_1/capacitor_5_2/buffer_digital_1/in clock_0/gnd 2.58f
C54 capacitors_5_1/capacitor_5_1/buffer_and_gate_0/and_gate_0/a_n78_396# clock_0/gnd 2.34f
C55 capacitors_5_1/capacitor_5_1/buffer_and_gate_0/buffer_0/a_1436_1552# clock_0/gnd 9.98f
C56 capacitors_5_1/capacitor_5_1/buffer_digital_1/in clock_0/gnd 2.58f
C57 capacitors_5_1/capacitor_5_0/buffer_and_gate_0/and_gate_0/a_n78_396# clock_0/gnd 2.34f
C58 capacitors_5_1/capacitor_5_0/buffer_and_gate_0/buffer_0/a_1436_1552# clock_0/gnd 9.98f
C59 capacitors_5_1/capacitor_5_0/buffer_digital_1/in clock_0/gnd 2.58f
C60 nmos_dnw3_0/out2 clock_0/gnd 16f
C61 capacitors_5_1/capacitor_5_7/buffer_and_gate_0/and_gate_0/a_n78_396# clock_0/gnd 2.34f
C62 clock_0/clk clock_0/gnd 86f
C63 clock_0/vdd clock_0/gnd 0.458p
C64 capacitors_5_1/capacitor_5_7/buffer_and_gate_0/buffer_0/a_1436_1552# clock_0/gnd 9.98f
C65 capacitors_5_1/capacitor_5_7/buffer_digital_1/in clock_0/gnd 2.58f
C66 capacitors_5_1/capacitor_5_6/buffer_and_gate_0/and_gate_0/a_n78_396# clock_0/gnd 2.34f
C67 capacitors_5_1/capacitor_5_6/buffer_and_gate_0/buffer_0/a_1436_1552# clock_0/gnd 9.98f
C68 capacitors_5_1/capacitor_5_6/buffer_digital_1/in clock_0/gnd 2.58f
C69 capacitors_5_1/capacitor_5_5/buffer_and_gate_0/and_gate_0/a_n78_396# clock_0/gnd 2.34f
C70 capacitors_5_1/capacitor_5_5/buffer_and_gate_0/buffer_0/a_1436_1552# clock_0/gnd 9.98f
C71 capacitors_5_1/capacitor_5_5/buffer_digital_1/in clock_0/gnd 2.58f
C72 nmos_dnw3_0/clk clock_0/gnd 2.53f
.ends

.subckt cp2_buffer2 buffer_digital_3/in charge_pump_reverse_0/capacitors_5_1/capacitor_5_1/i1
+ charge_pump_reverse_0/nmos_dnw3_0/vin charge_pump_reverse_0/capacitors_5_1/capacitor_5_2/i1
+ charge_pump_reverse_0/capacitors_5_1/capacitor_5_3/i1 charge_pump_reverse_0/capacitors_5_1/capacitor_5_4/i1
+ buffer_digital_3/VDD charge_pump_reverse_0/nmos_dnw3_0/vs charge_pump_reverse_0/m1_11946_n452#
+ charge_pump_reverse_0/capacitors_5_1/capacitor_5_5/i1 charge_pump_reverse_0/capacitors_5_1/capacitor_5_7/i1
+ buffer_digital_2/i charge_pump_reverse_0/capacitors_5_1/capacitor_5_0/i1 VSUBS charge_pump_reverse_0/capacitors_5_1/capacitor_5_6/i1
Xpmos_decap_10_10 VSUBS buffer_digital_3/VDD VSUBS pmos_decap_10
Xpmos_decap_10_11 VSUBS buffer_digital_3/VDD VSUBS pmos_decap_10
Xpmos_decap_10_12 VSUBS buffer_digital_3/VDD VSUBS pmos_decap_10
Xpmos_decap_10_13 VSUBS buffer_digital_3/VDD VSUBS pmos_decap_10
Xpmos_decap_10_14 VSUBS buffer_digital_3/VDD VSUBS pmos_decap_10
Xpmos_decap_10_15 VSUBS buffer_digital_3/VDD VSUBS pmos_decap_10
Xbuffer_digital_2 buffer_digital_2/i buffer_digital_3/i buffer_digital_3/VDD VSUBS
+ buffer_digital
Xbuffer_digital_3 buffer_digital_3/i buffer_digital_3/in buffer_digital_3/VDD VSUBS
+ buffer_digital
Xnmos_decap_10_0 buffer_digital_3/VDD VSUBS VSUBS nmos_decap_10
Xnmos_decap_10_1 buffer_digital_3/VDD VSUBS VSUBS nmos_decap_10
Xcharge_pump_reverse_0 charge_pump_reverse_0/m1_11946_n452# charge_pump_reverse_0/nmos_dnw3_0/vin
+ charge_pump_reverse_0/capacitors_5_1/capacitor_5_2/i1 charge_pump_reverse_0/capacitors_5_1/capacitor_5_3/i1
+ VSUBS charge_pump_reverse_0/capacitors_5_1/capacitor_5_4/i1 charge_pump_reverse_0/capacitors_5_1/capacitor_5_5/i1
+ buffer_digital_3/in buffer_digital_3/VDD charge_pump_reverse_0/capacitors_5_1/capacitor_5_0/i1
+ charge_pump_reverse_0/capacitors_5_1/capacitor_5_7/i1 VSUBS charge_pump_reverse_0/capacitors_5_1/capacitor_5_6/i1
+ charge_pump_reverse_0/capacitors_5_1/capacitor_5_1/i1 charge_pump_reverse_0/nmos_dnw3_0/vs
+ charge_pump_reverse
Xnmos_decap_10_2 buffer_digital_3/VDD VSUBS VSUBS nmos_decap_10
Xnmos_decap_10_3 buffer_digital_3/VDD VSUBS VSUBS nmos_decap_10
Xnmos_decap_10_4 buffer_digital_3/VDD VSUBS VSUBS nmos_decap_10
Xnmos_decap_10_5 buffer_digital_3/VDD VSUBS VSUBS nmos_decap_10
Xnmos_decap_10_6 buffer_digital_3/VDD VSUBS VSUBS nmos_decap_10
Xnmos_decap_10_7 buffer_digital_3/VDD VSUBS VSUBS nmos_decap_10
Xnmos_decap_10_8 buffer_digital_3/VDD VSUBS VSUBS nmos_decap_10
Xnmos_decap_10_9 buffer_digital_3/VDD VSUBS VSUBS nmos_decap_10
Xpmos_decap_10_0 VSUBS buffer_digital_3/VDD VSUBS pmos_decap_10
Xpmos_decap_10_1 VSUBS buffer_digital_3/VDD VSUBS pmos_decap_10
Xpmos_decap_10_2 VSUBS buffer_digital_3/VDD VSUBS pmos_decap_10
Xpmos_decap_10_3 VSUBS buffer_digital_3/VDD VSUBS pmos_decap_10
Xpmos_decap_10_4 VSUBS buffer_digital_3/VDD VSUBS pmos_decap_10
Xpmos_decap_10_5 VSUBS buffer_digital_3/VDD VSUBS pmos_decap_10
Xpmos_decap_10_6 VSUBS buffer_digital_3/VDD VSUBS pmos_decap_10
Xpmos_decap_10_7 VSUBS buffer_digital_3/VDD VSUBS pmos_decap_10
Xpmos_decap_10_9 VSUBS buffer_digital_3/VDD VSUBS pmos_decap_10
Xpmos_decap_10_8 VSUBS buffer_digital_3/VDD VSUBS pmos_decap_10
C0 charge_pump_reverse_0/clock_0/clkb buffer_digital_3/VDD 3.55f
C1 buffer_digital_3/VDD buffer_digital_3/in 5.15f
C2 buffer_digital_3/VDD buffer_digital_2/i 3.65f
C3 charge_pump_reverse_0/nmos_dnw3_0/vs VSUBS 18.8f
C4 charge_pump_reverse_0/clock_0/a_2432_n962# VSUBS 8.68f **FLOATING
C5 charge_pump_reverse_0/clock_0/a_2020_n482# VSUBS 2.57f **FLOATING
C6 charge_pump_reverse_0/clock_0/a_344_102# VSUBS 2.81f
C7 charge_pump_reverse_0/clock_0/a_2402_572# VSUBS 2.17f
C8 charge_pump_reverse_0/clock_0/a_344_n986# VSUBS 2.38f
C9 buffer_digital_3/in VSUBS 11.4f
C10 charge_pump_reverse_0/clock_0/a_3246_118# VSUBS 6.83f
C11 charge_pump_reverse_0/nmos_dnw3_0/vin VSUBS 2.46f
C12 charge_pump_reverse_0/nmos_dnw3_0/clkb VSUBS 2.23f
C13 charge_pump_reverse_0/capacitors_5_0/capacitor_5_4/buffer_and_gate_0/and_gate_0/a_n78_396# VSUBS 2.34f
C14 charge_pump_reverse_0/capacitors_5_0/capacitor_5_4/buffer_and_gate_0/buffer_0/a_1436_1552# VSUBS 9.98f
C15 charge_pump_reverse_0/capacitors_5_0/capacitor_5_4/buffer_digital_1/in VSUBS 2.58f
C16 charge_pump_reverse_0/capacitors_5_0/capacitor_5_3/buffer_and_gate_0/and_gate_0/a_n78_396# VSUBS 2.34f
C17 charge_pump_reverse_0/capacitors_5_0/capacitor_5_3/buffer_and_gate_0/buffer_0/a_1436_1552# VSUBS 9.98f
C18 charge_pump_reverse_0/capacitors_5_0/capacitor_5_3/buffer_digital_1/in VSUBS 2.58f
C19 charge_pump_reverse_0/capacitors_5_0/capacitor_5_2/buffer_and_gate_0/and_gate_0/a_n78_396# VSUBS 2.34f
C20 charge_pump_reverse_0/capacitors_5_0/capacitor_5_2/buffer_and_gate_0/buffer_0/a_1436_1552# VSUBS 9.98f
C21 charge_pump_reverse_0/capacitors_5_0/capacitor_5_2/buffer_digital_1/in VSUBS 2.58f
C22 charge_pump_reverse_0/capacitors_5_0/capacitor_5_1/buffer_and_gate_0/and_gate_0/a_n78_396# VSUBS 2.34f
C23 charge_pump_reverse_0/capacitors_5_0/capacitor_5_1/buffer_and_gate_0/buffer_0/a_1436_1552# VSUBS 9.98f
C24 charge_pump_reverse_0/capacitors_5_0/capacitor_5_1/buffer_digital_1/in VSUBS 2.58f
C25 charge_pump_reverse_0/capacitors_5_0/capacitor_5_0/buffer_and_gate_0/and_gate_0/a_n78_396# VSUBS 2.34f
C26 charge_pump_reverse_0/capacitors_5_0/capacitor_5_0/buffer_and_gate_0/buffer_0/a_1436_1552# VSUBS 9.98f
C27 charge_pump_reverse_0/capacitors_5_0/capacitor_5_0/buffer_digital_1/in VSUBS 2.58f
C28 charge_pump_reverse_0/nmos_dnw3_0/out1 VSUBS 15.1f
C29 charge_pump_reverse_0/capacitors_5_0/capacitor_5_7/buffer_and_gate_0/and_gate_0/a_n78_396# VSUBS 2.34f
C30 charge_pump_reverse_0/clock_0/clkb VSUBS 90.5f
C31 charge_pump_reverse_0/capacitors_5_0/capacitor_5_7/buffer_and_gate_0/buffer_0/a_1436_1552# VSUBS 9.98f
C32 charge_pump_reverse_0/capacitors_5_0/capacitor_5_7/buffer_digital_1/in VSUBS 2.58f
C33 charge_pump_reverse_0/capacitors_5_0/capacitor_5_6/buffer_and_gate_0/and_gate_0/a_n78_396# VSUBS 2.34f
C34 charge_pump_reverse_0/capacitors_5_0/capacitor_5_6/buffer_and_gate_0/buffer_0/a_1436_1552# VSUBS 9.98f
C35 charge_pump_reverse_0/capacitors_5_0/capacitor_5_6/buffer_digital_1/in VSUBS 2.58f
C36 charge_pump_reverse_0/capacitors_5_0/capacitor_5_5/buffer_and_gate_0/and_gate_0/a_n78_396# VSUBS 2.34f
C37 charge_pump_reverse_0/capacitors_5_0/capacitor_5_5/buffer_and_gate_0/buffer_0/a_1436_1552# VSUBS 9.98f
C38 charge_pump_reverse_0/capacitors_5_0/capacitor_5_5/buffer_digital_1/in VSUBS 2.58f
C39 charge_pump_reverse_0/capacitors_5_1/capacitor_5_4/buffer_and_gate_0/and_gate_0/a_n78_396# VSUBS 2.34f
C40 charge_pump_reverse_0/capacitors_5_1/capacitor_5_4/buffer_and_gate_0/buffer_0/a_1436_1552# VSUBS 9.98f
C41 charge_pump_reverse_0/capacitors_5_1/capacitor_5_4/buffer_digital_1/in VSUBS 2.58f
C42 charge_pump_reverse_0/capacitors_5_1/capacitor_5_3/buffer_and_gate_0/and_gate_0/a_n78_396# VSUBS 2.34f
C43 charge_pump_reverse_0/capacitors_5_1/capacitor_5_3/buffer_and_gate_0/buffer_0/a_1436_1552# VSUBS 9.98f
C44 charge_pump_reverse_0/capacitors_5_1/capacitor_5_3/buffer_digital_1/in VSUBS 2.58f
C45 charge_pump_reverse_0/capacitors_5_1/capacitor_5_2/buffer_and_gate_0/and_gate_0/a_n78_396# VSUBS 2.34f
C46 charge_pump_reverse_0/capacitors_5_1/capacitor_5_2/buffer_and_gate_0/buffer_0/a_1436_1552# VSUBS 9.98f
C47 charge_pump_reverse_0/capacitors_5_1/capacitor_5_2/buffer_digital_1/in VSUBS 2.58f
C48 charge_pump_reverse_0/capacitors_5_1/capacitor_5_1/buffer_and_gate_0/and_gate_0/a_n78_396# VSUBS 2.34f
C49 charge_pump_reverse_0/capacitors_5_1/capacitor_5_1/buffer_and_gate_0/buffer_0/a_1436_1552# VSUBS 9.98f
C50 charge_pump_reverse_0/capacitors_5_1/capacitor_5_1/buffer_digital_1/in VSUBS 2.58f
C51 charge_pump_reverse_0/capacitors_5_1/capacitor_5_0/buffer_and_gate_0/and_gate_0/a_n78_396# VSUBS 2.34f
C52 charge_pump_reverse_0/capacitors_5_1/capacitor_5_0/buffer_and_gate_0/buffer_0/a_1436_1552# VSUBS 9.98f
C53 charge_pump_reverse_0/capacitors_5_1/capacitor_5_0/buffer_digital_1/in VSUBS 2.58f
C54 charge_pump_reverse_0/nmos_dnw3_0/out2 VSUBS 14.8f
C55 charge_pump_reverse_0/capacitors_5_1/capacitor_5_7/buffer_and_gate_0/and_gate_0/a_n78_396# VSUBS 2.34f
C56 charge_pump_reverse_0/clock_0/clk VSUBS 84.6f
C57 buffer_digital_3/VDD VSUBS 0.547p
C58 charge_pump_reverse_0/capacitors_5_1/capacitor_5_7/buffer_and_gate_0/buffer_0/a_1436_1552# VSUBS 9.98f
C59 charge_pump_reverse_0/capacitors_5_1/capacitor_5_7/buffer_digital_1/in VSUBS 2.58f
C60 charge_pump_reverse_0/capacitors_5_1/capacitor_5_6/buffer_and_gate_0/and_gate_0/a_n78_396# VSUBS 2.34f
C61 charge_pump_reverse_0/capacitors_5_1/capacitor_5_6/buffer_and_gate_0/buffer_0/a_1436_1552# VSUBS 9.98f
C62 charge_pump_reverse_0/capacitors_5_1/capacitor_5_6/buffer_digital_1/in VSUBS 2.58f
C63 charge_pump_reverse_0/capacitors_5_1/capacitor_5_5/buffer_and_gate_0/and_gate_0/a_n78_396# VSUBS 2.34f
C64 charge_pump_reverse_0/capacitors_5_1/capacitor_5_5/buffer_and_gate_0/buffer_0/a_1436_1552# VSUBS 9.98f
C65 charge_pump_reverse_0/capacitors_5_1/capacitor_5_5/buffer_digital_1/in VSUBS 2.58f
C66 charge_pump_reverse_0/nmos_dnw3_0/clk VSUBS 2.43f
C67 buffer_digital_2/i VSUBS 10.7f
.ends

.subckt cp2_buffer_5stage cp2_buffer1_0/charge_pump_0/vin cp2_buffer1_1/charge_pump_0/vin
+ cp2_buffer1_1/charge_pump_0/out cp2_buffer1_2/charge_pump_0/in8 cp2_buffer1_2/charge_pump_0/in1
+ cp2_buffer1_2/charge_pump_0/vs cp2_buffer1_2/charge_pump_0/in2 cp2_buffer1_0/charge_pump_0/out
+ cp2_buffer1_2/charge_pump_0/in3 cp2_buffer2_0/charge_pump_reverse_0/nmos_dnw3_0/vs
+ cp2_buffer1_1/charge_pump_0/vs cp2_buffer2_1/charge_pump_reverse_0/nmos_dnw3_0/vs
+ cp2_buffer1_2/charge_pump_0/in4 cp2_buffer1_2/charge_pump_0/out cp2_buffer1_2/buffer_digital_0/in
+ cp2_buffer1_2/charge_pump_0/in5 cp2_buffer1_2/charge_pump_0/in7 cp2_buffer1_0/charge_pump_0/vs
+ cp2_buffer2_1/buffer_digital_3/VDD cp2_buffer1_2/charge_pump_0/in6 cp2_buffer1_0/buffer_digital_1/i
+ cp2_buffer1_2/charge_pump_0/a_18057_18271# VSUBS
Xcp2_buffer1_0 cp2_buffer1_0/charge_pump_0/a_18057_18271# cp2_buffer1_2/charge_pump_0/in4
+ cp2_buffer2_0/buffer_digital_2/i cp2_buffer1_2/charge_pump_0/in5 cp2_buffer1_0/charge_pump_0/vin
+ cp2_buffer1_0/charge_pump_0/out cp2_buffer1_2/charge_pump_0/in6 cp2_buffer1_2/charge_pump_0/in7
+ cp2_buffer1_0/charge_pump_0/vs cp2_buffer1_2/charge_pump_0/in8 cp2_buffer1_2/charge_pump_0/in1
+ cp2_buffer1_2/charge_pump_0/in3 cp2_buffer1_2/charge_pump_0/in2 cp2_buffer1_0/buffer_digital_1/i
+ VSUBS cp2_buffer2_1/buffer_digital_3/VDD cp2_buffer1
Xcp2_buffer1_1 cp2_buffer1_1/charge_pump_0/a_18057_18271# cp2_buffer1_2/charge_pump_0/in4
+ cp2_buffer2_1/buffer_digital_2/i cp2_buffer1_2/charge_pump_0/in5 cp2_buffer1_1/charge_pump_0/vin
+ cp2_buffer1_1/charge_pump_0/out cp2_buffer1_2/charge_pump_0/in6 cp2_buffer1_2/charge_pump_0/in7
+ cp2_buffer1_1/charge_pump_0/vs cp2_buffer1_2/charge_pump_0/in8 cp2_buffer1_2/charge_pump_0/in1
+ cp2_buffer1_2/charge_pump_0/in3 cp2_buffer1_2/charge_pump_0/in2 cp2_buffer1_1/buffer_digital_1/i
+ VSUBS cp2_buffer2_1/buffer_digital_3/VDD cp2_buffer1
Xcp2_buffer1_2 cp2_buffer1_2/charge_pump_0/a_18057_18271# cp2_buffer1_2/charge_pump_0/in4
+ cp2_buffer1_2/buffer_digital_0/in cp2_buffer1_2/charge_pump_0/in5 cp2_buffer1_2/charge_pump_0/vin
+ cp2_buffer1_2/charge_pump_0/out cp2_buffer1_2/charge_pump_0/in6 cp2_buffer1_2/charge_pump_0/in7
+ cp2_buffer1_2/charge_pump_0/vs cp2_buffer1_2/charge_pump_0/in8 cp2_buffer1_2/charge_pump_0/in1
+ cp2_buffer1_2/charge_pump_0/in3 cp2_buffer1_2/charge_pump_0/in2 cp2_buffer1_2/buffer_digital_1/i
+ VSUBS cp2_buffer2_1/buffer_digital_3/VDD cp2_buffer1
Xcp2_buffer2_0 cp2_buffer1_1/buffer_digital_1/i cp2_buffer1_2/charge_pump_0/in7 cp2_buffer1_0/charge_pump_0/out
+ cp2_buffer1_2/charge_pump_0/in6 cp2_buffer1_2/charge_pump_0/in5 cp2_buffer1_2/charge_pump_0/in4
+ cp2_buffer2_1/buffer_digital_3/VDD cp2_buffer2_0/charge_pump_reverse_0/nmos_dnw3_0/vs
+ cp2_buffer1_1/charge_pump_0/vin cp2_buffer1_2/charge_pump_0/in3 cp2_buffer1_2/charge_pump_0/in1
+ cp2_buffer2_0/buffer_digital_2/i cp2_buffer1_2/charge_pump_0/in8 VSUBS cp2_buffer1_2/charge_pump_0/in2
+ cp2_buffer2
Xcp2_buffer2_1 cp2_buffer1_2/buffer_digital_1/i cp2_buffer1_2/charge_pump_0/in7 cp2_buffer1_1/charge_pump_0/out
+ cp2_buffer1_2/charge_pump_0/in6 cp2_buffer1_2/charge_pump_0/in5 cp2_buffer1_2/charge_pump_0/in4
+ cp2_buffer2_1/buffer_digital_3/VDD cp2_buffer2_1/charge_pump_reverse_0/nmos_dnw3_0/vs
+ cp2_buffer1_2/charge_pump_0/vin cp2_buffer1_2/charge_pump_0/in3 cp2_buffer1_2/charge_pump_0/in1
+ cp2_buffer2_1/buffer_digital_2/i cp2_buffer1_2/charge_pump_0/in8 VSUBS cp2_buffer1_2/charge_pump_0/in2
+ cp2_buffer2
C0 cp2_buffer1_2/charge_pump_0/in8 cp2_buffer2_1/buffer_digital_3/VDD 4.65f
C1 cp2_buffer1_2/charge_pump_0/in1 cp2_buffer2_1/buffer_digital_3/VDD 4.32f
C2 cp2_buffer1_2/charge_pump_0/in2 cp2_buffer2_1/buffer_digital_3/VDD 4.4f
C3 cp2_buffer1_2/charge_pump_0/in3 cp2_buffer2_1/buffer_digital_3/VDD 4.42f
C4 cp2_buffer1_2/charge_pump_0/in7 cp2_buffer2_1/buffer_digital_3/VDD 4.45f
C5 cp2_buffer1_2/charge_pump_0/in4 cp2_buffer2_1/buffer_digital_3/VDD 4.39f
C6 cp2_buffer1_2/charge_pump_0/in5 cp2_buffer2_1/buffer_digital_3/VDD 4.39f
C7 cp2_buffer1_2/charge_pump_0/in6 cp2_buffer2_1/buffer_digital_3/VDD 4.45f
C8 cp2_buffer2_1/charge_pump_reverse_0/nmos_dnw3_0/vs cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 18.8f
C9 cp2_buffer2_1/charge_pump_reverse_0/clock_0/a_2432_n962# cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 8.68f **FLOATING
C10 cp2_buffer2_1/charge_pump_reverse_0/clock_0/a_2020_n482# cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.57f **FLOATING
C11 cp2_buffer2_1/charge_pump_reverse_0/clock_0/a_344_102# cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.81f
C12 cp2_buffer2_1/charge_pump_reverse_0/clock_0/a_2402_572# cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.17f
C13 cp2_buffer2_1/charge_pump_reverse_0/clock_0/a_344_n986# cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.38f
C14 cp2_buffer1_2/buffer_digital_1/i cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 8.96f
C15 cp2_buffer2_1/charge_pump_reverse_0/clock_0/a_3246_118# cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 6.83f
C16 cp2_buffer1_1/charge_pump_0/out cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 3.88f
C17 cp2_buffer2_1/charge_pump_reverse_0/nmos_dnw3_0/clkb cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.23f
C18 cp2_buffer2_1/charge_pump_reverse_0/capacitors_5_0/capacitor_5_4/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.34f
C19 cp2_buffer2_1/charge_pump_reverse_0/capacitors_5_0/capacitor_5_4/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.98f
C20 cp2_buffer2_1/charge_pump_reverse_0/capacitors_5_0/capacitor_5_4/buffer_digital_1/in cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.58f
C21 cp2_buffer2_1/charge_pump_reverse_0/capacitors_5_0/capacitor_5_3/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.34f
C22 cp2_buffer2_1/charge_pump_reverse_0/capacitors_5_0/capacitor_5_3/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.98f
C23 cp2_buffer2_1/charge_pump_reverse_0/capacitors_5_0/capacitor_5_3/buffer_digital_1/in cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.58f
C24 cp2_buffer2_1/charge_pump_reverse_0/capacitors_5_0/capacitor_5_2/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.34f
C25 cp2_buffer2_1/charge_pump_reverse_0/capacitors_5_0/capacitor_5_2/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.98f
C26 cp2_buffer2_1/charge_pump_reverse_0/capacitors_5_0/capacitor_5_2/buffer_digital_1/in cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.58f
C27 cp2_buffer2_1/charge_pump_reverse_0/capacitors_5_0/capacitor_5_1/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.34f
C28 cp2_buffer2_1/charge_pump_reverse_0/capacitors_5_0/capacitor_5_1/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.98f
C29 cp2_buffer2_1/charge_pump_reverse_0/capacitors_5_0/capacitor_5_1/buffer_digital_1/in cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.58f
C30 cp2_buffer2_1/charge_pump_reverse_0/capacitors_5_0/capacitor_5_0/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.34f
C31 cp2_buffer2_1/charge_pump_reverse_0/capacitors_5_0/capacitor_5_0/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.98f
C32 cp2_buffer2_1/charge_pump_reverse_0/capacitors_5_0/capacitor_5_0/buffer_digital_1/in cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.58f
C33 cp2_buffer2_1/charge_pump_reverse_0/nmos_dnw3_0/out1 cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 15.1f
C34 cp2_buffer2_1/charge_pump_reverse_0/capacitors_5_0/capacitor_5_7/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.34f
C35 cp2_buffer2_1/charge_pump_reverse_0/clock_0/clkb cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 91f
C36 cp2_buffer2_1/charge_pump_reverse_0/capacitors_5_0/capacitor_5_7/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.98f
C37 cp2_buffer2_1/charge_pump_reverse_0/capacitors_5_0/capacitor_5_7/buffer_digital_1/in cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.58f
C38 cp2_buffer2_1/charge_pump_reverse_0/capacitors_5_0/capacitor_5_6/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.34f
C39 cp2_buffer2_1/charge_pump_reverse_0/capacitors_5_0/capacitor_5_6/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.98f
C40 cp2_buffer2_1/charge_pump_reverse_0/capacitors_5_0/capacitor_5_6/buffer_digital_1/in cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.58f
C41 cp2_buffer2_1/charge_pump_reverse_0/capacitors_5_0/capacitor_5_5/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.34f
C42 cp2_buffer2_1/charge_pump_reverse_0/capacitors_5_0/capacitor_5_5/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.98f
C43 cp2_buffer2_1/charge_pump_reverse_0/capacitors_5_0/capacitor_5_5/buffer_digital_1/in cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.58f
C44 cp2_buffer2_1/charge_pump_reverse_0/capacitors_5_1/capacitor_5_4/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.34f
C45 cp2_buffer2_1/charge_pump_reverse_0/capacitors_5_1/capacitor_5_4/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.98f
C46 cp2_buffer2_1/charge_pump_reverse_0/capacitors_5_1/capacitor_5_4/buffer_digital_1/in cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.58f
C47 cp2_buffer2_1/charge_pump_reverse_0/capacitors_5_1/capacitor_5_3/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.34f
C48 cp2_buffer2_1/charge_pump_reverse_0/capacitors_5_1/capacitor_5_3/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.98f
C49 cp2_buffer2_1/charge_pump_reverse_0/capacitors_5_1/capacitor_5_3/buffer_digital_1/in cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.58f
C50 cp2_buffer2_1/charge_pump_reverse_0/capacitors_5_1/capacitor_5_2/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.34f
C51 cp2_buffer2_1/charge_pump_reverse_0/capacitors_5_1/capacitor_5_2/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.98f
C52 cp2_buffer2_1/charge_pump_reverse_0/capacitors_5_1/capacitor_5_2/buffer_digital_1/in cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.58f
C53 cp2_buffer2_1/charge_pump_reverse_0/capacitors_5_1/capacitor_5_1/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.34f
C54 cp2_buffer2_1/charge_pump_reverse_0/capacitors_5_1/capacitor_5_1/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.98f
C55 cp2_buffer2_1/charge_pump_reverse_0/capacitors_5_1/capacitor_5_1/buffer_digital_1/in cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.58f
C56 cp2_buffer2_1/charge_pump_reverse_0/capacitors_5_1/capacitor_5_0/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.34f
C57 cp2_buffer2_1/charge_pump_reverse_0/capacitors_5_1/capacitor_5_0/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.98f
C58 cp2_buffer2_1/charge_pump_reverse_0/capacitors_5_1/capacitor_5_0/buffer_digital_1/in cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.58f
C59 cp2_buffer2_1/charge_pump_reverse_0/nmos_dnw3_0/out2 cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 14.8f
C60 cp2_buffer2_1/charge_pump_reverse_0/capacitors_5_1/capacitor_5_7/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.34f
C61 cp2_buffer2_1/charge_pump_reverse_0/clock_0/clk cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 84.5f
C62 cp2_buffer2_1/charge_pump_reverse_0/capacitors_5_1/capacitor_5_7/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.98f
C63 cp2_buffer2_1/charge_pump_reverse_0/capacitors_5_1/capacitor_5_7/buffer_digital_1/in cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.58f
C64 cp2_buffer2_1/charge_pump_reverse_0/capacitors_5_1/capacitor_5_6/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.34f
C65 cp2_buffer2_1/charge_pump_reverse_0/capacitors_5_1/capacitor_5_6/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.98f
C66 cp2_buffer2_1/charge_pump_reverse_0/capacitors_5_1/capacitor_5_6/buffer_digital_1/in cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.58f
C67 cp2_buffer2_1/charge_pump_reverse_0/capacitors_5_1/capacitor_5_5/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.34f
C68 cp2_buffer2_1/charge_pump_reverse_0/capacitors_5_1/capacitor_5_5/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.98f
C69 cp2_buffer2_1/charge_pump_reverse_0/capacitors_5_1/capacitor_5_5/buffer_digital_1/in cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.58f
C70 cp2_buffer2_1/charge_pump_reverse_0/nmos_dnw3_0/clk cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.43f
C71 cp2_buffer2_0/charge_pump_reverse_0/nmos_dnw3_0/vs cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 18.8f
C72 cp2_buffer2_0/charge_pump_reverse_0/clock_0/a_2432_n962# cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 8.68f **FLOATING
C73 cp2_buffer2_0/charge_pump_reverse_0/clock_0/a_2020_n482# cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.57f **FLOATING
C74 cp2_buffer2_0/charge_pump_reverse_0/clock_0/a_344_102# cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.81f
C75 cp2_buffer2_0/charge_pump_reverse_0/clock_0/a_2402_572# cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.17f
C76 cp2_buffer2_0/charge_pump_reverse_0/clock_0/a_344_n986# cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.38f
C77 cp2_buffer1_1/buffer_digital_1/i cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 8.79f
C78 cp2_buffer2_0/charge_pump_reverse_0/clock_0/a_3246_118# cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 6.83f
C79 cp2_buffer1_0/charge_pump_0/out cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 4.36f
C80 cp2_buffer2_0/charge_pump_reverse_0/nmos_dnw3_0/clkb cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.23f
C81 cp2_buffer2_0/charge_pump_reverse_0/capacitors_5_0/capacitor_5_4/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.34f
C82 cp2_buffer2_0/charge_pump_reverse_0/capacitors_5_0/capacitor_5_4/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.98f
C83 cp2_buffer2_0/charge_pump_reverse_0/capacitors_5_0/capacitor_5_4/buffer_digital_1/in cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.58f
C84 cp2_buffer2_0/charge_pump_reverse_0/capacitors_5_0/capacitor_5_3/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.34f
C85 cp2_buffer2_0/charge_pump_reverse_0/capacitors_5_0/capacitor_5_3/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.98f
C86 cp2_buffer2_0/charge_pump_reverse_0/capacitors_5_0/capacitor_5_3/buffer_digital_1/in cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.58f
C87 cp2_buffer2_0/charge_pump_reverse_0/capacitors_5_0/capacitor_5_2/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.34f
C88 cp2_buffer2_0/charge_pump_reverse_0/capacitors_5_0/capacitor_5_2/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.98f
C89 cp2_buffer2_0/charge_pump_reverse_0/capacitors_5_0/capacitor_5_2/buffer_digital_1/in cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.58f
C90 cp2_buffer2_0/charge_pump_reverse_0/capacitors_5_0/capacitor_5_1/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.34f
C91 cp2_buffer2_0/charge_pump_reverse_0/capacitors_5_0/capacitor_5_1/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.98f
C92 cp2_buffer2_0/charge_pump_reverse_0/capacitors_5_0/capacitor_5_1/buffer_digital_1/in cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.58f
C93 cp2_buffer2_0/charge_pump_reverse_0/capacitors_5_0/capacitor_5_0/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.34f
C94 cp2_buffer2_0/charge_pump_reverse_0/capacitors_5_0/capacitor_5_0/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.98f
C95 cp2_buffer2_0/charge_pump_reverse_0/capacitors_5_0/capacitor_5_0/buffer_digital_1/in cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.58f
C96 cp2_buffer2_0/charge_pump_reverse_0/nmos_dnw3_0/out1 cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 15.1f
C97 cp2_buffer2_0/charge_pump_reverse_0/capacitors_5_0/capacitor_5_7/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.34f
C98 cp2_buffer2_0/charge_pump_reverse_0/clock_0/clkb cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 90.9f
C99 cp2_buffer2_0/charge_pump_reverse_0/capacitors_5_0/capacitor_5_7/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.98f
C100 cp2_buffer2_0/charge_pump_reverse_0/capacitors_5_0/capacitor_5_7/buffer_digital_1/in cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.58f
C101 cp2_buffer2_0/charge_pump_reverse_0/capacitors_5_0/capacitor_5_6/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.34f
C102 cp2_buffer2_0/charge_pump_reverse_0/capacitors_5_0/capacitor_5_6/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.98f
C103 cp2_buffer2_0/charge_pump_reverse_0/capacitors_5_0/capacitor_5_6/buffer_digital_1/in cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.58f
C104 cp2_buffer2_0/charge_pump_reverse_0/capacitors_5_0/capacitor_5_5/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.34f
C105 cp2_buffer2_0/charge_pump_reverse_0/capacitors_5_0/capacitor_5_5/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.98f
C106 cp2_buffer2_0/charge_pump_reverse_0/capacitors_5_0/capacitor_5_5/buffer_digital_1/in cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.58f
C107 cp2_buffer1_2/charge_pump_0/in3 cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 14.7f
C108 cp2_buffer2_0/charge_pump_reverse_0/capacitors_5_1/capacitor_5_4/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.34f
C109 cp2_buffer2_0/charge_pump_reverse_0/capacitors_5_1/capacitor_5_4/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.98f
C110 cp2_buffer2_0/charge_pump_reverse_0/capacitors_5_1/capacitor_5_4/buffer_digital_1/in cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.58f
C111 cp2_buffer2_0/charge_pump_reverse_0/capacitors_5_1/capacitor_5_3/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.34f
C112 cp2_buffer2_0/charge_pump_reverse_0/capacitors_5_1/capacitor_5_3/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.98f
C113 cp2_buffer2_0/charge_pump_reverse_0/capacitors_5_1/capacitor_5_3/buffer_digital_1/in cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.58f
C114 cp2_buffer2_0/charge_pump_reverse_0/capacitors_5_1/capacitor_5_2/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.34f
C115 cp2_buffer2_0/charge_pump_reverse_0/capacitors_5_1/capacitor_5_2/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.98f
C116 cp2_buffer2_0/charge_pump_reverse_0/capacitors_5_1/capacitor_5_2/buffer_digital_1/in cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.58f
C117 cp2_buffer2_0/charge_pump_reverse_0/capacitors_5_1/capacitor_5_1/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.34f
C118 cp2_buffer2_0/charge_pump_reverse_0/capacitors_5_1/capacitor_5_1/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.98f
C119 cp2_buffer2_0/charge_pump_reverse_0/capacitors_5_1/capacitor_5_1/buffer_digital_1/in cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.58f
C120 cp2_buffer2_0/charge_pump_reverse_0/capacitors_5_1/capacitor_5_0/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.34f
C121 cp2_buffer2_0/charge_pump_reverse_0/capacitors_5_1/capacitor_5_0/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.98f
C122 cp2_buffer2_0/charge_pump_reverse_0/capacitors_5_1/capacitor_5_0/buffer_digital_1/in cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.58f
C123 cp2_buffer1_2/charge_pump_0/in8 cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 14.2f
C124 cp2_buffer2_0/charge_pump_reverse_0/nmos_dnw3_0/out2 cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 14.8f
C125 cp2_buffer2_0/charge_pump_reverse_0/capacitors_5_1/capacitor_5_7/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.34f
C126 cp2_buffer2_0/charge_pump_reverse_0/clock_0/clk cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 84.6f
C127 cp2_buffer2_0/charge_pump_reverse_0/capacitors_5_1/capacitor_5_7/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.98f
C128 cp2_buffer2_0/charge_pump_reverse_0/capacitors_5_1/capacitor_5_7/buffer_digital_1/in cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.58f
C129 cp2_buffer2_0/charge_pump_reverse_0/capacitors_5_1/capacitor_5_6/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.34f
C130 cp2_buffer2_0/charge_pump_reverse_0/capacitors_5_1/capacitor_5_6/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.98f
C131 cp2_buffer2_0/charge_pump_reverse_0/capacitors_5_1/capacitor_5_6/buffer_digital_1/in cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.58f
C132 cp2_buffer2_0/charge_pump_reverse_0/capacitors_5_1/capacitor_5_5/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.34f
C133 cp2_buffer2_0/charge_pump_reverse_0/capacitors_5_1/capacitor_5_5/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.98f
C134 cp2_buffer2_0/charge_pump_reverse_0/capacitors_5_1/capacitor_5_5/buffer_digital_1/in cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.58f
C135 cp2_buffer2_0/charge_pump_reverse_0/nmos_dnw3_0/clk cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.43f
C136 cp2_buffer1_2/charge_pump_0/vin cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 3.49f
C137 cp2_buffer1_2/charge_pump_0/vs cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 19f
C138 cp2_buffer1_2/charge_pump_0/clock_0/a_2432_n962# cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 8.68f **FLOATING
C139 cp2_buffer1_2/charge_pump_0/clock_0/a_2020_n482# cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.57f **FLOATING
C140 cp2_buffer1_2/charge_pump_0/clock_0/a_344_102# cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.81f
C141 cp2_buffer1_2/charge_pump_0/clock_0/a_2402_572# cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.17f
C142 cp2_buffer1_2/charge_pump_0/clock_0/a_344_n986# cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.38f
C143 cp2_buffer1_2/buffer_digital_0/in cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 4.6f
C144 cp2_buffer1_2/charge_pump_0/clock_0/a_3246_118# cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 6.83f
C145 cp2_buffer1_2/charge_pump_0/g2 cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.44f
C146 cp2_buffer1_2/charge_pump_0/capacitors_5_0/capacitor_5_4/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.34f
C147 cp2_buffer1_2/charge_pump_0/capacitors_5_0/capacitor_5_4/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.98f
C148 cp2_buffer1_2/charge_pump_0/capacitors_5_0/capacitor_5_4/buffer_digital_1/in cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.58f
C149 cp2_buffer1_2/charge_pump_0/capacitors_5_0/capacitor_5_3/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.34f
C150 cp2_buffer1_2/charge_pump_0/capacitors_5_0/capacitor_5_3/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.98f
C151 cp2_buffer1_2/charge_pump_0/capacitors_5_0/capacitor_5_3/buffer_digital_1/in cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.58f
C152 cp2_buffer1_2/charge_pump_0/capacitors_5_0/capacitor_5_2/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.34f
C153 cp2_buffer1_2/charge_pump_0/capacitors_5_0/capacitor_5_2/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.98f
C154 cp2_buffer1_2/charge_pump_0/capacitors_5_0/capacitor_5_2/buffer_digital_1/in cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.58f
C155 cp2_buffer1_2/charge_pump_0/capacitors_5_0/capacitor_5_1/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.34f
C156 cp2_buffer1_2/charge_pump_0/capacitors_5_0/capacitor_5_1/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.98f
C157 cp2_buffer1_2/charge_pump_0/capacitors_5_0/capacitor_5_1/buffer_digital_1/in cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.58f
C158 cp2_buffer1_2/charge_pump_0/capacitors_5_0/capacitor_5_0/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.34f
C159 cp2_buffer1_2/charge_pump_0/capacitors_5_0/capacitor_5_0/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.98f
C160 cp2_buffer1_2/charge_pump_0/capacitors_5_0/capacitor_5_0/buffer_digital_1/in cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.58f
C161 cp2_buffer1_2/charge_pump_0/input1 cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 15f
C162 cp2_buffer1_2/charge_pump_0/capacitors_5_0/capacitor_5_7/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.34f
C163 cp2_buffer1_2/charge_pump_0/clk cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 82.5f
C164 cp2_buffer1_2/charge_pump_0/capacitors_5_0/capacitor_5_7/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.98f
C165 cp2_buffer1_2/charge_pump_0/capacitors_5_0/capacitor_5_7/buffer_digital_1/in cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.58f
C166 cp2_buffer1_2/charge_pump_0/capacitors_5_0/capacitor_5_6/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.34f
C167 cp2_buffer1_2/charge_pump_0/capacitors_5_0/capacitor_5_6/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.98f
C168 cp2_buffer1_2/charge_pump_0/capacitors_5_0/capacitor_5_6/buffer_digital_1/in cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.58f
C169 cp2_buffer1_2/charge_pump_0/in7 cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 14.8f
C170 cp2_buffer1_2/charge_pump_0/capacitors_5_0/capacitor_5_5/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.34f
C171 cp2_buffer1_2/charge_pump_0/capacitors_5_0/capacitor_5_5/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.98f
C172 cp2_buffer1_2/charge_pump_0/capacitors_5_0/capacitor_5_5/buffer_digital_1/in cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.58f
C173 cp2_buffer1_2/charge_pump_0/capacitors_5_1/capacitor_5_4/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.34f
C174 cp2_buffer1_2/charge_pump_0/capacitors_5_1/capacitor_5_4/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.98f
C175 cp2_buffer1_2/charge_pump_0/capacitors_5_1/capacitor_5_4/buffer_digital_1/in cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.58f
C176 cp2_buffer1_2/charge_pump_0/capacitors_5_1/capacitor_5_3/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.34f
C177 cp2_buffer1_2/charge_pump_0/capacitors_5_1/capacitor_5_3/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.98f
C178 cp2_buffer1_2/charge_pump_0/capacitors_5_1/capacitor_5_3/buffer_digital_1/in cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.58f
C179 cp2_buffer1_2/charge_pump_0/capacitors_5_1/capacitor_5_2/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.34f
C180 cp2_buffer1_2/charge_pump_0/capacitors_5_1/capacitor_5_2/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.98f
C181 cp2_buffer1_2/charge_pump_0/capacitors_5_1/capacitor_5_2/buffer_digital_1/in cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.58f
C182 cp2_buffer1_2/charge_pump_0/capacitors_5_1/capacitor_5_1/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.34f
C183 cp2_buffer1_2/charge_pump_0/capacitors_5_1/capacitor_5_1/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.98f
C184 cp2_buffer1_2/charge_pump_0/capacitors_5_1/capacitor_5_1/buffer_digital_1/in cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.58f
C185 cp2_buffer1_2/charge_pump_0/capacitors_5_1/capacitor_5_0/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.34f
C186 cp2_buffer1_2/charge_pump_0/capacitors_5_1/capacitor_5_0/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.98f
C187 cp2_buffer1_2/charge_pump_0/capacitors_5_1/capacitor_5_0/buffer_digital_1/in cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.58f
C188 cp2_buffer1_2/charge_pump_0/input2 cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 14.4f
C189 cp2_buffer1_2/charge_pump_0/capacitors_5_1/capacitor_5_7/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.34f
C190 cp2_buffer1_2/charge_pump_0/clkb cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 83.8f
C191 cp2_buffer1_2/charge_pump_0/capacitors_5_1/capacitor_5_7/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.98f
C192 cp2_buffer1_2/charge_pump_0/capacitors_5_1/capacitor_5_7/buffer_digital_1/in cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.58f
C193 cp2_buffer1_2/charge_pump_0/capacitors_5_1/capacitor_5_6/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.34f
C194 cp2_buffer1_2/charge_pump_0/capacitors_5_1/capacitor_5_6/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.98f
C195 cp2_buffer1_2/charge_pump_0/capacitors_5_1/capacitor_5_6/buffer_digital_1/in cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.58f
C196 cp2_buffer1_2/charge_pump_0/capacitors_5_1/capacitor_5_5/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.34f
C197 cp2_buffer1_2/charge_pump_0/capacitors_5_1/capacitor_5_5/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.98f
C198 cp2_buffer1_2/charge_pump_0/capacitors_5_1/capacitor_5_5/buffer_digital_1/in cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.58f
C199 cp2_buffer1_2/charge_pump_0/g1 cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.63f
C200 cp2_buffer1_1/charge_pump_0/vin cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 3.62f
C201 cp2_buffer1_1/charge_pump_0/vs cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 19f
C202 cp2_buffer1_1/charge_pump_0/clock_0/a_2432_n962# cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 8.68f **FLOATING
C203 cp2_buffer1_1/charge_pump_0/clock_0/a_2020_n482# cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.57f **FLOATING
C204 cp2_buffer1_1/charge_pump_0/clock_0/a_344_102# cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.81f
C205 cp2_buffer1_1/charge_pump_0/clock_0/a_2402_572# cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.17f
C206 cp2_buffer1_1/charge_pump_0/clock_0/a_344_n986# cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.38f
C207 cp2_buffer2_1/buffer_digital_2/i cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 7.16f
C208 cp2_buffer1_1/charge_pump_0/clock_0/a_3246_118# cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 6.83f
C209 cp2_buffer1_1/charge_pump_0/g2 cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.44f
C210 cp2_buffer1_1/charge_pump_0/capacitors_5_0/capacitor_5_4/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.34f
C211 cp2_buffer1_1/charge_pump_0/capacitors_5_0/capacitor_5_4/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.98f
C212 cp2_buffer1_1/charge_pump_0/capacitors_5_0/capacitor_5_4/buffer_digital_1/in cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.58f
C213 cp2_buffer1_2/charge_pump_0/in5 cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 14.7f
C214 cp2_buffer1_1/charge_pump_0/capacitors_5_0/capacitor_5_3/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.34f
C215 cp2_buffer1_1/charge_pump_0/capacitors_5_0/capacitor_5_3/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.98f
C216 cp2_buffer1_1/charge_pump_0/capacitors_5_0/capacitor_5_3/buffer_digital_1/in cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.58f
C217 cp2_buffer1_1/charge_pump_0/capacitors_5_0/capacitor_5_2/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.34f
C218 cp2_buffer1_1/charge_pump_0/capacitors_5_0/capacitor_5_2/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.98f
C219 cp2_buffer1_1/charge_pump_0/capacitors_5_0/capacitor_5_2/buffer_digital_1/in cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.58f
C220 cp2_buffer1_1/charge_pump_0/capacitors_5_0/capacitor_5_1/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.34f
C221 cp2_buffer1_1/charge_pump_0/capacitors_5_0/capacitor_5_1/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.98f
C222 cp2_buffer1_1/charge_pump_0/capacitors_5_0/capacitor_5_1/buffer_digital_1/in cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.58f
C223 cp2_buffer1_2/charge_pump_0/in2 cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 14.8f
C224 cp2_buffer1_1/charge_pump_0/capacitors_5_0/capacitor_5_0/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.34f
C225 cp2_buffer1_1/charge_pump_0/capacitors_5_0/capacitor_5_0/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.98f
C226 cp2_buffer1_1/charge_pump_0/capacitors_5_0/capacitor_5_0/buffer_digital_1/in cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.58f
C227 cp2_buffer1_1/charge_pump_0/input1 cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 15f
C228 cp2_buffer1_1/charge_pump_0/capacitors_5_0/capacitor_5_7/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.34f
C229 cp2_buffer1_1/charge_pump_0/clk cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 82.5f
C230 cp2_buffer1_1/charge_pump_0/capacitors_5_0/capacitor_5_7/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.98f
C231 cp2_buffer1_1/charge_pump_0/capacitors_5_0/capacitor_5_7/buffer_digital_1/in cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.58f
C232 cp2_buffer1_1/charge_pump_0/capacitors_5_0/capacitor_5_6/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.34f
C233 cp2_buffer1_1/charge_pump_0/capacitors_5_0/capacitor_5_6/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.98f
C234 cp2_buffer1_1/charge_pump_0/capacitors_5_0/capacitor_5_6/buffer_digital_1/in cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.58f
C235 cp2_buffer1_1/charge_pump_0/capacitors_5_0/capacitor_5_5/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.34f
C236 cp2_buffer1_1/charge_pump_0/capacitors_5_0/capacitor_5_5/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.98f
C237 cp2_buffer1_1/charge_pump_0/capacitors_5_0/capacitor_5_5/buffer_digital_1/in cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.58f
C238 cp2_buffer1_2/charge_pump_0/in6 cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 14.7f
C239 cp2_buffer1_1/charge_pump_0/capacitors_5_1/capacitor_5_4/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.34f
C240 cp2_buffer1_1/charge_pump_0/capacitors_5_1/capacitor_5_4/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.98f
C241 cp2_buffer1_1/charge_pump_0/capacitors_5_1/capacitor_5_4/buffer_digital_1/in cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.58f
C242 cp2_buffer1_1/charge_pump_0/capacitors_5_1/capacitor_5_3/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.34f
C243 cp2_buffer1_1/charge_pump_0/capacitors_5_1/capacitor_5_3/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.98f
C244 cp2_buffer1_1/charge_pump_0/capacitors_5_1/capacitor_5_3/buffer_digital_1/in cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.58f
C245 cp2_buffer1_1/charge_pump_0/capacitors_5_1/capacitor_5_2/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.34f
C246 cp2_buffer1_1/charge_pump_0/capacitors_5_1/capacitor_5_2/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.98f
C247 cp2_buffer1_1/charge_pump_0/capacitors_5_1/capacitor_5_2/buffer_digital_1/in cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.58f
C248 cp2_buffer1_1/charge_pump_0/capacitors_5_1/capacitor_5_1/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.34f
C249 cp2_buffer1_1/charge_pump_0/capacitors_5_1/capacitor_5_1/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.98f
C250 cp2_buffer1_1/charge_pump_0/capacitors_5_1/capacitor_5_1/buffer_digital_1/in cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.58f
C251 cp2_buffer1_1/charge_pump_0/capacitors_5_1/capacitor_5_0/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.34f
C252 cp2_buffer1_1/charge_pump_0/capacitors_5_1/capacitor_5_0/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.98f
C253 cp2_buffer1_1/charge_pump_0/capacitors_5_1/capacitor_5_0/buffer_digital_1/in cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.58f
C254 cp2_buffer1_1/charge_pump_0/input2 cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 14.4f
C255 cp2_buffer1_1/charge_pump_0/capacitors_5_1/capacitor_5_7/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.34f
C256 cp2_buffer1_1/charge_pump_0/clkb cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 83.9f
C257 cp2_buffer1_1/charge_pump_0/capacitors_5_1/capacitor_5_7/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.98f
C258 cp2_buffer1_1/charge_pump_0/capacitors_5_1/capacitor_5_7/buffer_digital_1/in cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.58f
C259 cp2_buffer1_1/charge_pump_0/capacitors_5_1/capacitor_5_6/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.34f
C260 cp2_buffer1_1/charge_pump_0/capacitors_5_1/capacitor_5_6/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.98f
C261 cp2_buffer1_1/charge_pump_0/capacitors_5_1/capacitor_5_6/buffer_digital_1/in cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.58f
C262 cp2_buffer1_1/charge_pump_0/capacitors_5_1/capacitor_5_5/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.34f
C263 cp2_buffer1_1/charge_pump_0/capacitors_5_1/capacitor_5_5/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.98f
C264 cp2_buffer1_1/charge_pump_0/capacitors_5_1/capacitor_5_5/buffer_digital_1/in cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.58f
C265 cp2_buffer1_1/charge_pump_0/g1 cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.63f
C266 cp2_buffer1_0/buffer_digital_1/i cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 4.02f
C267 cp2_buffer1_0/charge_pump_0/vs cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 19f
C268 cp2_buffer1_0/charge_pump_0/clock_0/a_2432_n962# cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 8.68f **FLOATING
C269 cp2_buffer1_0/charge_pump_0/clock_0/a_2020_n482# cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.57f **FLOATING
C270 cp2_buffer1_0/charge_pump_0/clock_0/a_344_102# cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.81f
C271 cp2_buffer1_0/charge_pump_0/clock_0/a_2402_572# cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.17f
C272 cp2_buffer1_0/charge_pump_0/clock_0/a_344_n986# cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.38f
C273 cp2_buffer2_0/buffer_digital_2/i cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 8.22f
C274 cp2_buffer1_0/charge_pump_0/clock_0/a_3246_118# cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 6.83f
C275 cp2_buffer1_0/charge_pump_0/g2 cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.44f
C276 cp2_buffer1_0/charge_pump_0/capacitors_5_0/capacitor_5_4/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.34f
C277 cp2_buffer1_0/charge_pump_0/capacitors_5_0/capacitor_5_4/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.98f
C278 cp2_buffer1_0/charge_pump_0/capacitors_5_0/capacitor_5_4/buffer_digital_1/in cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.58f
C279 cp2_buffer1_0/charge_pump_0/capacitors_5_0/capacitor_5_3/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.34f
C280 cp2_buffer1_0/charge_pump_0/capacitors_5_0/capacitor_5_3/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.98f
C281 cp2_buffer1_0/charge_pump_0/capacitors_5_0/capacitor_5_3/buffer_digital_1/in cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.58f
C282 cp2_buffer1_2/charge_pump_0/in4 cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 14.7f
C283 cp2_buffer1_0/charge_pump_0/capacitors_5_0/capacitor_5_2/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.34f
C284 cp2_buffer1_0/charge_pump_0/capacitors_5_0/capacitor_5_2/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.98f
C285 cp2_buffer1_0/charge_pump_0/capacitors_5_0/capacitor_5_2/buffer_digital_1/in cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.58f
C286 cp2_buffer1_0/charge_pump_0/capacitors_5_0/capacitor_5_1/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.34f
C287 cp2_buffer1_0/charge_pump_0/capacitors_5_0/capacitor_5_1/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.98f
C288 cp2_buffer1_0/charge_pump_0/capacitors_5_0/capacitor_5_1/buffer_digital_1/in cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.58f
C289 cp2_buffer1_0/charge_pump_0/capacitors_5_0/capacitor_5_0/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.34f
C290 cp2_buffer1_0/charge_pump_0/capacitors_5_0/capacitor_5_0/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.98f
C291 cp2_buffer1_0/charge_pump_0/capacitors_5_0/capacitor_5_0/buffer_digital_1/in cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.58f
C292 cp2_buffer1_2/charge_pump_0/in1 cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 14.1f
C293 cp2_buffer1_0/charge_pump_0/input1 cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 15f
C294 cp2_buffer1_0/charge_pump_0/capacitors_5_0/capacitor_5_7/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.34f
C295 cp2_buffer1_0/charge_pump_0/clk cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 82.1f
C296 cp2_buffer2_1/buffer_digital_3/VDD cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.56p
C297 cp2_buffer1_0/charge_pump_0/capacitors_5_0/capacitor_5_7/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.99f
C298 cp2_buffer1_0/charge_pump_0/capacitors_5_0/capacitor_5_7/buffer_digital_1/in cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.58f
C299 cp2_buffer1_0/charge_pump_0/capacitors_5_0/capacitor_5_6/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.34f
C300 cp2_buffer1_0/charge_pump_0/capacitors_5_0/capacitor_5_6/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.98f
C301 cp2_buffer1_0/charge_pump_0/capacitors_5_0/capacitor_5_6/buffer_digital_1/in cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.58f
C302 cp2_buffer1_0/charge_pump_0/capacitors_5_0/capacitor_5_5/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.34f
C303 cp2_buffer1_0/charge_pump_0/capacitors_5_0/capacitor_5_5/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.98f
C304 cp2_buffer1_0/charge_pump_0/capacitors_5_0/capacitor_5_5/buffer_digital_1/in cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.58f
C305 cp2_buffer1_0/charge_pump_0/capacitors_5_1/capacitor_5_4/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.34f
C306 cp2_buffer1_0/charge_pump_0/capacitors_5_1/capacitor_5_4/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.98f
C307 cp2_buffer1_0/charge_pump_0/capacitors_5_1/capacitor_5_4/buffer_digital_1/in cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.58f
C308 cp2_buffer1_0/charge_pump_0/capacitors_5_1/capacitor_5_3/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.34f
C309 cp2_buffer1_0/charge_pump_0/capacitors_5_1/capacitor_5_3/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.98f
C310 cp2_buffer1_0/charge_pump_0/capacitors_5_1/capacitor_5_3/buffer_digital_1/in cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.58f
C311 cp2_buffer1_0/charge_pump_0/capacitors_5_1/capacitor_5_2/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.34f
C312 cp2_buffer1_0/charge_pump_0/capacitors_5_1/capacitor_5_2/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.98f
C313 cp2_buffer1_0/charge_pump_0/capacitors_5_1/capacitor_5_2/buffer_digital_1/in cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.58f
C314 cp2_buffer1_0/charge_pump_0/capacitors_5_1/capacitor_5_1/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.34f
C315 cp2_buffer1_0/charge_pump_0/capacitors_5_1/capacitor_5_1/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.98f
C316 cp2_buffer1_0/charge_pump_0/capacitors_5_1/capacitor_5_1/buffer_digital_1/in cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.58f
C317 cp2_buffer1_0/charge_pump_0/capacitors_5_1/capacitor_5_0/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.34f
C318 cp2_buffer1_0/charge_pump_0/capacitors_5_1/capacitor_5_0/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.98f
C319 cp2_buffer1_0/charge_pump_0/capacitors_5_1/capacitor_5_0/buffer_digital_1/in cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.58f
C320 cp2_buffer1_0/charge_pump_0/input2 cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 14.4f
C321 cp2_buffer1_0/charge_pump_0/capacitors_5_1/capacitor_5_7/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.34f
C322 cp2_buffer1_0/charge_pump_0/clkb cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 83.9f
C323 cp2_buffer1_0/charge_pump_0/capacitors_5_1/capacitor_5_7/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.98f
C324 cp2_buffer1_0/charge_pump_0/capacitors_5_1/capacitor_5_7/buffer_digital_1/in cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.58f
C325 cp2_buffer1_0/charge_pump_0/capacitors_5_1/capacitor_5_6/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.34f
C326 cp2_buffer1_0/charge_pump_0/capacitors_5_1/capacitor_5_6/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.98f
C327 cp2_buffer1_0/charge_pump_0/capacitors_5_1/capacitor_5_6/buffer_digital_1/in cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.58f
C328 cp2_buffer1_0/charge_pump_0/capacitors_5_1/capacitor_5_5/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.34f
C329 cp2_buffer1_0/charge_pump_0/capacitors_5_1/capacitor_5_5/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.98f
C330 cp2_buffer1_0/charge_pump_0/capacitors_5_1/capacitor_5_5/buffer_digital_1/in cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.58f
C331 cp2_buffer1_0/charge_pump_0/g1 cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.63f
.ends

.subckt reconfigurable_CP
Xscanchain_0 scanchain_0/data_out[0] scanchain_0/data_out[1] scanchain_0/data_out[2]
+ scanchain_0/data_out[3] scanchain_0/data_out[4] scanchain_0/data_out[5] scanchain_0/data_out[6]
+ scanchain_0/data_out[7] scanchain_0/scan_out scanchain_0/VDD VSUBS scanchain
Xcp1_buffer_5stage_0 scanchain_0/data_out[1] scanchain_0/data_out[7] scanchain_0/data_out[6]
+ scanchain_0/data_out[5] scanchain_0/data_out[0] scanchain_0/data_out[4] cp2_buffer_5stage_0/cp2_buffer1_0/charge_pump_0/vin
+ cp1_buffer_5stage_0/cp1_buffer1_reverse_1/charge_pump1_reverse_0/nmos_dnw3_0/vs
+ cp1_buffer_5stage_0/cp1_buffer1_0/clk_in scanchain_0/data_out[3] cp1_buffer_5stage_0/cp1_buffer1_reverse_0/charge_pump1_reverse_0/nmos_dnw3_0/vs
+ cp1_buffer_5stage_0/cp1_buffer1_0/charge_pump1_0/vin cp1_buffer_5stage_0/cp1_buffer1_1/charge_pump1_0/vin
+ scanchain_0/VDD VSUBS scanchain_0/data_out[2] cp2_buffer_5stage_0/cp2_buffer1_0/charge_pump_0/vs
+ cp1_buffer_5stage
Xcp2_buffer_5stage_0 cp2_buffer_5stage_0/cp2_buffer1_0/charge_pump_0/vin cp2_buffer_5stage_0/cp2_buffer1_1/charge_pump_0/vin
+ cp2_buffer_5stage_1/cp2_buffer1_0/charge_pump_0/vs scanchain_0/data_out[0] scanchain_0/data_out[7]
+ cp2_buffer_5stage_1/cp2_buffer1_0/charge_pump_0/vs scanchain_0/data_out[6] cp2_buffer_5stage_0/cp2_buffer1_1/charge_pump_0/vs
+ scanchain_0/data_out[5] cp2_buffer_5stage_0/cp2_buffer1_0/charge_pump_0/vin cp2_buffer_5stage_0/cp2_buffer1_1/charge_pump_0/vs
+ cp2_buffer_5stage_0/cp2_buffer1_1/charge_pump_0/vin scanchain_0/data_out[4] cp2_buffer_5stage_1/cp2_buffer1_0/charge_pump_0/vin
+ cp2_buffer_5stage_0/cp2_buffer1_2/buffer_digital_0/in scanchain_0/data_out[3] scanchain_0/data_out[1]
+ cp2_buffer_5stage_0/cp2_buffer1_0/charge_pump_0/vs scanchain_0/VDD scanchain_0/data_out[2]
+ cp2_buffer_5stage_0/cp2_buffer1_0/buffer_digital_1/i cp2_buffer_5stage_0/cp2_buffer1_2/charge_pump_0/a_18057_18271#
+ VSUBS cp2_buffer_5stage
Xcp2_buffer_5stage_1 cp2_buffer_5stage_1/cp2_buffer1_0/charge_pump_0/vin cp2_buffer_5stage_1/cp2_buffer1_1/charge_pump_0/vin
+ cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/vs scanchain_0/data_out[7] scanchain_0/data_out[0]
+ cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/vs scanchain_0/data_out[1] cp2_buffer_5stage_1/cp2_buffer1_1/charge_pump_0/vs
+ scanchain_0/data_out[2] cp2_buffer_5stage_1/cp2_buffer1_0/charge_pump_0/vin cp2_buffer_5stage_1/cp2_buffer1_1/charge_pump_0/vs
+ cp2_buffer_5stage_1/cp2_buffer1_1/charge_pump_0/vin scanchain_0/data_out[3] cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/out
+ cp2_buffer_5stage_0/cp2_buffer1_0/buffer_digital_1/i scanchain_0/data_out[4] scanchain_0/data_out[6]
+ cp2_buffer_5stage_1/cp2_buffer1_0/charge_pump_0/vs scanchain_0/VDD scanchain_0/data_out[5]
+ cp1_buffer_5stage_0/cp1_buffer1_0/clk_in VSUBS VSUBS cp2_buffer_5stage
C0 scanchain_0/data_out[0] scanchain_0/data_out[7] 3.24f
C1 scanchain_0/data_out[4] scanchain_0/VDD 3.05f
C2 scanchain_0/data_out[0] scanchain_0/data_out[1] 13.4f
C3 scanchain_0/data_out[6] scanchain_0/data_out[2] 2.24f
C4 scanchain_0/VDD scanchain_0/data_out[7] 3.17f
C5 scanchain_0/data_out[6] scanchain_0/data_out[5] 8.2f
C6 scanchain_0/VDD scanchain_0/data_out[3] 2.63f
C7 scanchain_0/VDD scanchain_0/data_out[1] 2.86f
C8 scanchain_0/data_out[4] scanchain_0/data_out[3] 10.5f
C9 scanchain_0/VDD scanchain_0/data_out[2] 2.54f
C10 scanchain_0/data_out[6] scanchain_0/VDD 3.75f
C11 scanchain_0/VDD scanchain_0/data_out[5] 3.3f
C12 scanchain_0/VDD cp2_buffer_5stage_0/cp2_buffer1_0/buffer_digital_1/i 8.53f
C13 scanchain_0/data_out[4] scanchain_0/data_out[5] 9.18f
C14 cp1_buffer_5stage_0/cp1_buffer1_0/clk_in scanchain_0/VDD 9.99f
C15 scanchain_0/data_out[6] scanchain_0/data_out[7] 5.47f
C16 scanchain_0/data_out[0] scanchain_0/VDD 3.19f
C17 scanchain_0/data_out[3] scanchain_0/data_out[2] 9.12f
C18 scanchain_0/data_out[1] scanchain_0/data_out[2] 8.23f
C19 scanchain_0/data_out[6] scanchain_0/data_out[1] 2.69f
C20 cp2_buffer_5stage_1/cp2_buffer1_1/charge_pump_0/vin cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 23.5f
C21 cp2_buffer_5stage_1/cp2_buffer2_1/charge_pump_reverse_0/clock_0/a_2432_n962# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 8.68f **FLOATING
C22 cp2_buffer_5stage_1/cp2_buffer2_1/charge_pump_reverse_0/clock_0/a_2020_n482# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.57f **FLOATING
C23 cp2_buffer_5stage_1/cp2_buffer2_1/charge_pump_reverse_0/clock_0/a_344_102# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.81f
C24 cp2_buffer_5stage_1/cp2_buffer2_1/charge_pump_reverse_0/clock_0/a_2402_572# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.17f
C25 cp2_buffer_5stage_1/cp2_buffer2_1/charge_pump_reverse_0/clock_0/a_344_n986# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.38f
C26 cp2_buffer_5stage_1/cp2_buffer1_2/buffer_digital_1/i cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 7.41f
C27 cp2_buffer_5stage_1/cp2_buffer2_1/charge_pump_reverse_0/clock_0/a_3246_118# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 6.83f
C28 cp2_buffer_5stage_1/cp2_buffer2_1/charge_pump_reverse_0/nmos_dnw3_0/clkb cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.23f
C29 cp2_buffer_5stage_1/cp2_buffer2_1/charge_pump_reverse_0/capacitors_5_0/capacitor_5_4/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.34f
C30 cp2_buffer_5stage_1/cp2_buffer2_1/charge_pump_reverse_0/capacitors_5_0/capacitor_5_4/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.98f
C31 cp2_buffer_5stage_1/cp2_buffer2_1/charge_pump_reverse_0/capacitors_5_0/capacitor_5_4/buffer_digital_1/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.58f
C32 cp2_buffer_5stage_1/cp2_buffer2_1/charge_pump_reverse_0/capacitors_5_0/capacitor_5_3/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.34f
C33 cp2_buffer_5stage_1/cp2_buffer2_1/charge_pump_reverse_0/capacitors_5_0/capacitor_5_3/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.98f
C34 cp2_buffer_5stage_1/cp2_buffer2_1/charge_pump_reverse_0/capacitors_5_0/capacitor_5_3/buffer_digital_1/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.58f
C35 cp2_buffer_5stage_1/cp2_buffer2_1/charge_pump_reverse_0/capacitors_5_0/capacitor_5_2/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.34f
C36 cp2_buffer_5stage_1/cp2_buffer2_1/charge_pump_reverse_0/capacitors_5_0/capacitor_5_2/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.98f
C37 cp2_buffer_5stage_1/cp2_buffer2_1/charge_pump_reverse_0/capacitors_5_0/capacitor_5_2/buffer_digital_1/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.58f
C38 cp2_buffer_5stage_1/cp2_buffer2_1/charge_pump_reverse_0/capacitors_5_0/capacitor_5_1/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.34f
C39 cp2_buffer_5stage_1/cp2_buffer2_1/charge_pump_reverse_0/capacitors_5_0/capacitor_5_1/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.98f
C40 cp2_buffer_5stage_1/cp2_buffer2_1/charge_pump_reverse_0/capacitors_5_0/capacitor_5_1/buffer_digital_1/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.58f
C41 cp2_buffer_5stage_1/cp2_buffer2_1/charge_pump_reverse_0/capacitors_5_0/capacitor_5_0/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.34f
C42 cp2_buffer_5stage_1/cp2_buffer2_1/charge_pump_reverse_0/capacitors_5_0/capacitor_5_0/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.98f
C43 cp2_buffer_5stage_1/cp2_buffer2_1/charge_pump_reverse_0/capacitors_5_0/capacitor_5_0/buffer_digital_1/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.58f
C44 cp2_buffer_5stage_1/cp2_buffer2_1/charge_pump_reverse_0/nmos_dnw3_0/out1 cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 15.1f
C45 cp2_buffer_5stage_1/cp2_buffer2_1/charge_pump_reverse_0/capacitors_5_0/capacitor_5_7/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.34f
C46 cp2_buffer_5stage_1/cp2_buffer2_1/charge_pump_reverse_0/clock_0/clkb cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 90.9f
C47 cp2_buffer_5stage_1/cp2_buffer2_1/charge_pump_reverse_0/capacitors_5_0/capacitor_5_7/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.98f
C48 cp2_buffer_5stage_1/cp2_buffer2_1/charge_pump_reverse_0/capacitors_5_0/capacitor_5_7/buffer_digital_1/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.58f
C49 cp2_buffer_5stage_1/cp2_buffer2_1/charge_pump_reverse_0/capacitors_5_0/capacitor_5_6/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.34f
C50 cp2_buffer_5stage_1/cp2_buffer2_1/charge_pump_reverse_0/capacitors_5_0/capacitor_5_6/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.98f
C51 cp2_buffer_5stage_1/cp2_buffer2_1/charge_pump_reverse_0/capacitors_5_0/capacitor_5_6/buffer_digital_1/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.58f
C52 cp2_buffer_5stage_1/cp2_buffer2_1/charge_pump_reverse_0/capacitors_5_0/capacitor_5_5/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.34f
C53 cp2_buffer_5stage_1/cp2_buffer2_1/charge_pump_reverse_0/capacitors_5_0/capacitor_5_5/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.98f
C54 cp2_buffer_5stage_1/cp2_buffer2_1/charge_pump_reverse_0/capacitors_5_0/capacitor_5_5/buffer_digital_1/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.58f
C55 cp2_buffer_5stage_1/cp2_buffer2_1/charge_pump_reverse_0/capacitors_5_1/capacitor_5_4/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.34f
C56 cp2_buffer_5stage_1/cp2_buffer2_1/charge_pump_reverse_0/capacitors_5_1/capacitor_5_4/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.98f
C57 cp2_buffer_5stage_1/cp2_buffer2_1/charge_pump_reverse_0/capacitors_5_1/capacitor_5_4/buffer_digital_1/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.58f
C58 cp2_buffer_5stage_1/cp2_buffer2_1/charge_pump_reverse_0/capacitors_5_1/capacitor_5_3/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.34f
C59 cp2_buffer_5stage_1/cp2_buffer2_1/charge_pump_reverse_0/capacitors_5_1/capacitor_5_3/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.98f
C60 cp2_buffer_5stage_1/cp2_buffer2_1/charge_pump_reverse_0/capacitors_5_1/capacitor_5_3/buffer_digital_1/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.58f
C61 cp2_buffer_5stage_1/cp2_buffer2_1/charge_pump_reverse_0/capacitors_5_1/capacitor_5_2/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.34f
C62 cp2_buffer_5stage_1/cp2_buffer2_1/charge_pump_reverse_0/capacitors_5_1/capacitor_5_2/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.98f
C63 cp2_buffer_5stage_1/cp2_buffer2_1/charge_pump_reverse_0/capacitors_5_1/capacitor_5_2/buffer_digital_1/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.58f
C64 cp2_buffer_5stage_1/cp2_buffer2_1/charge_pump_reverse_0/capacitors_5_1/capacitor_5_1/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.34f
C65 cp2_buffer_5stage_1/cp2_buffer2_1/charge_pump_reverse_0/capacitors_5_1/capacitor_5_1/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.98f
C66 cp2_buffer_5stage_1/cp2_buffer2_1/charge_pump_reverse_0/capacitors_5_1/capacitor_5_1/buffer_digital_1/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.58f
C67 cp2_buffer_5stage_1/cp2_buffer2_1/charge_pump_reverse_0/capacitors_5_1/capacitor_5_0/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.34f
C68 cp2_buffer_5stage_1/cp2_buffer2_1/charge_pump_reverse_0/capacitors_5_1/capacitor_5_0/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.98f
C69 cp2_buffer_5stage_1/cp2_buffer2_1/charge_pump_reverse_0/capacitors_5_1/capacitor_5_0/buffer_digital_1/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.58f
C70 cp2_buffer_5stage_1/cp2_buffer2_1/charge_pump_reverse_0/nmos_dnw3_0/out2 cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 14.8f
C71 cp2_buffer_5stage_1/cp2_buffer2_1/charge_pump_reverse_0/capacitors_5_1/capacitor_5_7/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.34f
C72 cp2_buffer_5stage_1/cp2_buffer2_1/charge_pump_reverse_0/clock_0/clk cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 84.5f
C73 cp2_buffer_5stage_1/cp2_buffer2_1/charge_pump_reverse_0/capacitors_5_1/capacitor_5_7/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.98f
C74 cp2_buffer_5stage_1/cp2_buffer2_1/charge_pump_reverse_0/capacitors_5_1/capacitor_5_7/buffer_digital_1/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.58f
C75 cp2_buffer_5stage_1/cp2_buffer2_1/charge_pump_reverse_0/capacitors_5_1/capacitor_5_6/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.34f
C76 cp2_buffer_5stage_1/cp2_buffer2_1/charge_pump_reverse_0/capacitors_5_1/capacitor_5_6/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.98f
C77 cp2_buffer_5stage_1/cp2_buffer2_1/charge_pump_reverse_0/capacitors_5_1/capacitor_5_6/buffer_digital_1/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.58f
C78 cp2_buffer_5stage_1/cp2_buffer2_1/charge_pump_reverse_0/capacitors_5_1/capacitor_5_5/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.34f
C79 cp2_buffer_5stage_1/cp2_buffer2_1/charge_pump_reverse_0/capacitors_5_1/capacitor_5_5/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.98f
C80 cp2_buffer_5stage_1/cp2_buffer2_1/charge_pump_reverse_0/capacitors_5_1/capacitor_5_5/buffer_digital_1/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.58f
C81 cp2_buffer_5stage_1/cp2_buffer2_1/charge_pump_reverse_0/nmos_dnw3_0/clk cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.43f
C82 cp2_buffer_5stage_1/cp2_buffer1_0/charge_pump_0/vin cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 29.2f
C83 cp2_buffer_5stage_1/cp2_buffer2_0/charge_pump_reverse_0/clock_0/a_2432_n962# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 8.68f **FLOATING
C84 cp2_buffer_5stage_1/cp2_buffer2_0/charge_pump_reverse_0/clock_0/a_2020_n482# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.57f **FLOATING
C85 cp2_buffer_5stage_1/cp2_buffer2_0/charge_pump_reverse_0/clock_0/a_344_102# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.81f
C86 cp2_buffer_5stage_1/cp2_buffer2_0/charge_pump_reverse_0/clock_0/a_2402_572# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.17f
C87 cp2_buffer_5stage_1/cp2_buffer2_0/charge_pump_reverse_0/clock_0/a_344_n986# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.38f
C88 cp2_buffer_5stage_1/cp2_buffer1_1/buffer_digital_1/i cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 7.27f
C89 cp2_buffer_5stage_1/cp2_buffer2_0/charge_pump_reverse_0/clock_0/a_3246_118# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 6.83f
C90 cp2_buffer_5stage_1/cp2_buffer2_0/charge_pump_reverse_0/nmos_dnw3_0/clkb cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.23f
C91 cp2_buffer_5stage_1/cp2_buffer2_0/charge_pump_reverse_0/capacitors_5_0/capacitor_5_4/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.34f
C92 cp2_buffer_5stage_1/cp2_buffer2_0/charge_pump_reverse_0/capacitors_5_0/capacitor_5_4/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.98f
C93 cp2_buffer_5stage_1/cp2_buffer2_0/charge_pump_reverse_0/capacitors_5_0/capacitor_5_4/buffer_digital_1/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.58f
C94 cp2_buffer_5stage_1/cp2_buffer2_0/charge_pump_reverse_0/capacitors_5_0/capacitor_5_3/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.34f
C95 cp2_buffer_5stage_1/cp2_buffer2_0/charge_pump_reverse_0/capacitors_5_0/capacitor_5_3/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.98f
C96 cp2_buffer_5stage_1/cp2_buffer2_0/charge_pump_reverse_0/capacitors_5_0/capacitor_5_3/buffer_digital_1/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.58f
C97 cp2_buffer_5stage_1/cp2_buffer2_0/charge_pump_reverse_0/capacitors_5_0/capacitor_5_2/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.34f
C98 cp2_buffer_5stage_1/cp2_buffer2_0/charge_pump_reverse_0/capacitors_5_0/capacitor_5_2/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.98f
C99 cp2_buffer_5stage_1/cp2_buffer2_0/charge_pump_reverse_0/capacitors_5_0/capacitor_5_2/buffer_digital_1/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.58f
C100 cp2_buffer_5stage_1/cp2_buffer2_0/charge_pump_reverse_0/capacitors_5_0/capacitor_5_1/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.34f
C101 cp2_buffer_5stage_1/cp2_buffer2_0/charge_pump_reverse_0/capacitors_5_0/capacitor_5_1/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.98f
C102 cp2_buffer_5stage_1/cp2_buffer2_0/charge_pump_reverse_0/capacitors_5_0/capacitor_5_1/buffer_digital_1/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.58f
C103 cp2_buffer_5stage_1/cp2_buffer2_0/charge_pump_reverse_0/capacitors_5_0/capacitor_5_0/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.34f
C104 cp2_buffer_5stage_1/cp2_buffer2_0/charge_pump_reverse_0/capacitors_5_0/capacitor_5_0/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.98f
C105 cp2_buffer_5stage_1/cp2_buffer2_0/charge_pump_reverse_0/capacitors_5_0/capacitor_5_0/buffer_digital_1/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.58f
C106 cp2_buffer_5stage_1/cp2_buffer2_0/charge_pump_reverse_0/nmos_dnw3_0/out1 cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 15.1f
C107 cp2_buffer_5stage_1/cp2_buffer2_0/charge_pump_reverse_0/capacitors_5_0/capacitor_5_7/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.34f
C108 cp2_buffer_5stage_1/cp2_buffer2_0/charge_pump_reverse_0/clock_0/clkb cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 90.9f
C109 cp2_buffer_5stage_1/cp2_buffer2_0/charge_pump_reverse_0/capacitors_5_0/capacitor_5_7/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.98f
C110 cp2_buffer_5stage_1/cp2_buffer2_0/charge_pump_reverse_0/capacitors_5_0/capacitor_5_7/buffer_digital_1/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.58f
C111 cp2_buffer_5stage_1/cp2_buffer2_0/charge_pump_reverse_0/capacitors_5_0/capacitor_5_6/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.34f
C112 cp2_buffer_5stage_1/cp2_buffer2_0/charge_pump_reverse_0/capacitors_5_0/capacitor_5_6/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.98f
C113 cp2_buffer_5stage_1/cp2_buffer2_0/charge_pump_reverse_0/capacitors_5_0/capacitor_5_6/buffer_digital_1/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.58f
C114 cp2_buffer_5stage_1/cp2_buffer2_0/charge_pump_reverse_0/capacitors_5_0/capacitor_5_5/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.34f
C115 cp2_buffer_5stage_1/cp2_buffer2_0/charge_pump_reverse_0/capacitors_5_0/capacitor_5_5/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.98f
C116 cp2_buffer_5stage_1/cp2_buffer2_0/charge_pump_reverse_0/capacitors_5_0/capacitor_5_5/buffer_digital_1/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.58f
C117 scanchain_0/data_out[2] cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 38.9f
C118 cp2_buffer_5stage_1/cp2_buffer2_0/charge_pump_reverse_0/capacitors_5_1/capacitor_5_4/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.34f
C119 cp2_buffer_5stage_1/cp2_buffer2_0/charge_pump_reverse_0/capacitors_5_1/capacitor_5_4/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.98f
C120 cp2_buffer_5stage_1/cp2_buffer2_0/charge_pump_reverse_0/capacitors_5_1/capacitor_5_4/buffer_digital_1/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.58f
C121 cp2_buffer_5stage_1/cp2_buffer2_0/charge_pump_reverse_0/capacitors_5_1/capacitor_5_3/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.34f
C122 cp2_buffer_5stage_1/cp2_buffer2_0/charge_pump_reverse_0/capacitors_5_1/capacitor_5_3/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.98f
C123 cp2_buffer_5stage_1/cp2_buffer2_0/charge_pump_reverse_0/capacitors_5_1/capacitor_5_3/buffer_digital_1/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.58f
C124 cp2_buffer_5stage_1/cp2_buffer2_0/charge_pump_reverse_0/capacitors_5_1/capacitor_5_2/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.34f
C125 cp2_buffer_5stage_1/cp2_buffer2_0/charge_pump_reverse_0/capacitors_5_1/capacitor_5_2/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.98f
C126 cp2_buffer_5stage_1/cp2_buffer2_0/charge_pump_reverse_0/capacitors_5_1/capacitor_5_2/buffer_digital_1/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.58f
C127 cp2_buffer_5stage_1/cp2_buffer2_0/charge_pump_reverse_0/capacitors_5_1/capacitor_5_1/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.34f
C128 cp2_buffer_5stage_1/cp2_buffer2_0/charge_pump_reverse_0/capacitors_5_1/capacitor_5_1/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.98f
C129 cp2_buffer_5stage_1/cp2_buffer2_0/charge_pump_reverse_0/capacitors_5_1/capacitor_5_1/buffer_digital_1/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.58f
C130 cp2_buffer_5stage_1/cp2_buffer2_0/charge_pump_reverse_0/capacitors_5_1/capacitor_5_0/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.34f
C131 cp2_buffer_5stage_1/cp2_buffer2_0/charge_pump_reverse_0/capacitors_5_1/capacitor_5_0/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.98f
C132 cp2_buffer_5stage_1/cp2_buffer2_0/charge_pump_reverse_0/capacitors_5_1/capacitor_5_0/buffer_digital_1/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.58f
C133 scanchain_0/data_out[7] cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 54.1f
C134 cp2_buffer_5stage_1/cp2_buffer2_0/charge_pump_reverse_0/nmos_dnw3_0/out2 cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 14.8f
C135 cp2_buffer_5stage_1/cp2_buffer2_0/charge_pump_reverse_0/capacitors_5_1/capacitor_5_7/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.34f
C136 cp2_buffer_5stage_1/cp2_buffer2_0/charge_pump_reverse_0/clock_0/clk cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 84.5f
C137 cp2_buffer_5stage_1/cp2_buffer2_0/charge_pump_reverse_0/capacitors_5_1/capacitor_5_7/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.98f
C138 cp2_buffer_5stage_1/cp2_buffer2_0/charge_pump_reverse_0/capacitors_5_1/capacitor_5_7/buffer_digital_1/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.58f
C139 cp2_buffer_5stage_1/cp2_buffer2_0/charge_pump_reverse_0/capacitors_5_1/capacitor_5_6/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.34f
C140 cp2_buffer_5stage_1/cp2_buffer2_0/charge_pump_reverse_0/capacitors_5_1/capacitor_5_6/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.98f
C141 cp2_buffer_5stage_1/cp2_buffer2_0/charge_pump_reverse_0/capacitors_5_1/capacitor_5_6/buffer_digital_1/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.58f
C142 cp2_buffer_5stage_1/cp2_buffer2_0/charge_pump_reverse_0/capacitors_5_1/capacitor_5_5/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.34f
C143 cp2_buffer_5stage_1/cp2_buffer2_0/charge_pump_reverse_0/capacitors_5_1/capacitor_5_5/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.98f
C144 cp2_buffer_5stage_1/cp2_buffer2_0/charge_pump_reverse_0/capacitors_5_1/capacitor_5_5/buffer_digital_1/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.58f
C145 cp2_buffer_5stage_1/cp2_buffer2_0/charge_pump_reverse_0/nmos_dnw3_0/clk cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.43f
C146 cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/vin cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 3.28f
C147 cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/vs cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 23.7f
C148 cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/clock_0/a_2432_n962# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 8.68f **FLOATING
C149 cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/clock_0/a_2020_n482# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.57f **FLOATING
C150 cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/clock_0/a_344_102# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.81f
C151 cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/clock_0/a_2402_572# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.17f
C152 cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/clock_0/a_344_n986# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.38f
C153 cp2_buffer_5stage_0/cp2_buffer1_0/buffer_digital_1/i cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 11.4f
C154 cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/clock_0/a_3246_118# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 6.83f
C155 cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/g2 cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.44f
C156 cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/capacitors_5_0/capacitor_5_4/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.34f
C157 cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/capacitors_5_0/capacitor_5_4/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.98f
C158 cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/capacitors_5_0/capacitor_5_4/buffer_digital_1/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.58f
C159 cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/capacitors_5_0/capacitor_5_3/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.34f
C160 cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/capacitors_5_0/capacitor_5_3/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.98f
C161 cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/capacitors_5_0/capacitor_5_3/buffer_digital_1/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.58f
C162 cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/capacitors_5_0/capacitor_5_2/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.34f
C163 cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/capacitors_5_0/capacitor_5_2/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.98f
C164 cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/capacitors_5_0/capacitor_5_2/buffer_digital_1/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.58f
C165 cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/capacitors_5_0/capacitor_5_1/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.34f
C166 cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/capacitors_5_0/capacitor_5_1/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.98f
C167 cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/capacitors_5_0/capacitor_5_1/buffer_digital_1/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.58f
C168 cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/capacitors_5_0/capacitor_5_0/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.34f
C169 cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/capacitors_5_0/capacitor_5_0/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.98f
C170 cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/capacitors_5_0/capacitor_5_0/buffer_digital_1/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.58f
C171 cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/input1 cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 15f
C172 cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/capacitors_5_0/capacitor_5_7/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.34f
C173 cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/clk cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 82.3f
C174 cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/capacitors_5_0/capacitor_5_7/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.98f
C175 cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/capacitors_5_0/capacitor_5_7/buffer_digital_1/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.58f
C176 cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/capacitors_5_0/capacitor_5_6/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.34f
C177 cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/capacitors_5_0/capacitor_5_6/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.98f
C178 cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/capacitors_5_0/capacitor_5_6/buffer_digital_1/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.58f
C179 cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/capacitors_5_0/capacitor_5_5/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.34f
C180 cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/capacitors_5_0/capacitor_5_5/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.98f
C181 cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/capacitors_5_0/capacitor_5_5/buffer_digital_1/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.58f
C182 cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/capacitors_5_1/capacitor_5_4/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.34f
C183 cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/capacitors_5_1/capacitor_5_4/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.98f
C184 cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/capacitors_5_1/capacitor_5_4/buffer_digital_1/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.58f
C185 cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/capacitors_5_1/capacitor_5_3/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.34f
C186 cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/capacitors_5_1/capacitor_5_3/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.98f
C187 cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/capacitors_5_1/capacitor_5_3/buffer_digital_1/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.58f
C188 cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/capacitors_5_1/capacitor_5_2/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.34f
C189 cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/capacitors_5_1/capacitor_5_2/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.98f
C190 cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/capacitors_5_1/capacitor_5_2/buffer_digital_1/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.58f
C191 cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/capacitors_5_1/capacitor_5_1/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.34f
C192 cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/capacitors_5_1/capacitor_5_1/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.98f
C193 cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/capacitors_5_1/capacitor_5_1/buffer_digital_1/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.58f
C194 cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/capacitors_5_1/capacitor_5_0/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.34f
C195 cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/capacitors_5_1/capacitor_5_0/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.98f
C196 cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/capacitors_5_1/capacitor_5_0/buffer_digital_1/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.58f
C197 cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/input2 cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 14.4f
C198 cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/capacitors_5_1/capacitor_5_7/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.34f
C199 cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/clkb cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 83.9f
C200 cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/capacitors_5_1/capacitor_5_7/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.98f
C201 cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/capacitors_5_1/capacitor_5_7/buffer_digital_1/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.58f
C202 cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/capacitors_5_1/capacitor_5_6/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.34f
C203 cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/capacitors_5_1/capacitor_5_6/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.98f
C204 cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/capacitors_5_1/capacitor_5_6/buffer_digital_1/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.58f
C205 cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/capacitors_5_1/capacitor_5_5/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.34f
C206 cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/capacitors_5_1/capacitor_5_5/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.98f
C207 cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/capacitors_5_1/capacitor_5_5/buffer_digital_1/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.58f
C208 cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/g1 cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.63f
C209 cp2_buffer_5stage_1/cp2_buffer1_1/charge_pump_0/vs cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 24.1f
C210 cp2_buffer_5stage_1/cp2_buffer1_1/charge_pump_0/clock_0/a_2432_n962# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 8.68f **FLOATING
C211 cp2_buffer_5stage_1/cp2_buffer1_1/charge_pump_0/clock_0/a_2020_n482# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.57f **FLOATING
C212 cp2_buffer_5stage_1/cp2_buffer1_1/charge_pump_0/clock_0/a_344_102# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.81f
C213 cp2_buffer_5stage_1/cp2_buffer1_1/charge_pump_0/clock_0/a_2402_572# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.17f
C214 cp2_buffer_5stage_1/cp2_buffer1_1/charge_pump_0/clock_0/a_344_n986# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.38f
C215 cp2_buffer_5stage_1/cp2_buffer2_1/buffer_digital_2/i cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 6.84f
C216 cp2_buffer_5stage_1/cp2_buffer1_1/charge_pump_0/clock_0/a_3246_118# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 6.83f
C217 cp2_buffer_5stage_1/cp2_buffer1_1/charge_pump_0/g2 cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.44f
C218 cp2_buffer_5stage_1/cp2_buffer1_1/charge_pump_0/capacitors_5_0/capacitor_5_4/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.34f
C219 cp2_buffer_5stage_1/cp2_buffer1_1/charge_pump_0/capacitors_5_0/capacitor_5_4/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.98f
C220 cp2_buffer_5stage_1/cp2_buffer1_1/charge_pump_0/capacitors_5_0/capacitor_5_4/buffer_digital_1/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.58f
C221 cp2_buffer_5stage_1/cp2_buffer1_1/charge_pump_0/capacitors_5_0/capacitor_5_3/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.34f
C222 cp2_buffer_5stage_1/cp2_buffer1_1/charge_pump_0/capacitors_5_0/capacitor_5_3/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.98f
C223 cp2_buffer_5stage_1/cp2_buffer1_1/charge_pump_0/capacitors_5_0/capacitor_5_3/buffer_digital_1/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.58f
C224 cp2_buffer_5stage_1/cp2_buffer1_1/charge_pump_0/capacitors_5_0/capacitor_5_2/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.34f
C225 cp2_buffer_5stage_1/cp2_buffer1_1/charge_pump_0/capacitors_5_0/capacitor_5_2/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.98f
C226 cp2_buffer_5stage_1/cp2_buffer1_1/charge_pump_0/capacitors_5_0/capacitor_5_2/buffer_digital_1/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.58f
C227 cp2_buffer_5stage_1/cp2_buffer1_1/charge_pump_0/capacitors_5_0/capacitor_5_1/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.34f
C228 cp2_buffer_5stage_1/cp2_buffer1_1/charge_pump_0/capacitors_5_0/capacitor_5_1/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.98f
C229 cp2_buffer_5stage_1/cp2_buffer1_1/charge_pump_0/capacitors_5_0/capacitor_5_1/buffer_digital_1/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.58f
C230 scanchain_0/data_out[1] cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 36.9f
C231 cp2_buffer_5stage_1/cp2_buffer1_1/charge_pump_0/capacitors_5_0/capacitor_5_0/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.34f
C232 cp2_buffer_5stage_1/cp2_buffer1_1/charge_pump_0/capacitors_5_0/capacitor_5_0/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.98f
C233 cp2_buffer_5stage_1/cp2_buffer1_1/charge_pump_0/capacitors_5_0/capacitor_5_0/buffer_digital_1/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.58f
C234 cp2_buffer_5stage_1/cp2_buffer1_1/charge_pump_0/input1 cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 15f
C235 cp2_buffer_5stage_1/cp2_buffer1_1/charge_pump_0/capacitors_5_0/capacitor_5_7/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.34f
C236 cp2_buffer_5stage_1/cp2_buffer1_1/charge_pump_0/clk cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 82.3f
C237 cp2_buffer_5stage_1/cp2_buffer1_1/charge_pump_0/capacitors_5_0/capacitor_5_7/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.98f
C238 cp2_buffer_5stage_1/cp2_buffer1_1/charge_pump_0/capacitors_5_0/capacitor_5_7/buffer_digital_1/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.58f
C239 cp2_buffer_5stage_1/cp2_buffer1_1/charge_pump_0/capacitors_5_0/capacitor_5_6/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.34f
C240 cp2_buffer_5stage_1/cp2_buffer1_1/charge_pump_0/capacitors_5_0/capacitor_5_6/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.98f
C241 cp2_buffer_5stage_1/cp2_buffer1_1/charge_pump_0/capacitors_5_0/capacitor_5_6/buffer_digital_1/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.58f
C242 cp2_buffer_5stage_1/cp2_buffer1_1/charge_pump_0/capacitors_5_0/capacitor_5_5/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.34f
C243 cp2_buffer_5stage_1/cp2_buffer1_1/charge_pump_0/capacitors_5_0/capacitor_5_5/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.98f
C244 cp2_buffer_5stage_1/cp2_buffer1_1/charge_pump_0/capacitors_5_0/capacitor_5_5/buffer_digital_1/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.58f
C245 scanchain_0/data_out[5] cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 32.6f
C246 cp2_buffer_5stage_1/cp2_buffer1_1/charge_pump_0/capacitors_5_1/capacitor_5_4/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.34f
C247 cp2_buffer_5stage_1/cp2_buffer1_1/charge_pump_0/capacitors_5_1/capacitor_5_4/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.98f
C248 cp2_buffer_5stage_1/cp2_buffer1_1/charge_pump_0/capacitors_5_1/capacitor_5_4/buffer_digital_1/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.58f
C249 cp2_buffer_5stage_1/cp2_buffer1_1/charge_pump_0/capacitors_5_1/capacitor_5_3/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.34f
C250 cp2_buffer_5stage_1/cp2_buffer1_1/charge_pump_0/capacitors_5_1/capacitor_5_3/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.98f
C251 cp2_buffer_5stage_1/cp2_buffer1_1/charge_pump_0/capacitors_5_1/capacitor_5_3/buffer_digital_1/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.58f
C252 cp2_buffer_5stage_1/cp2_buffer1_1/charge_pump_0/capacitors_5_1/capacitor_5_2/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.34f
C253 cp2_buffer_5stage_1/cp2_buffer1_1/charge_pump_0/capacitors_5_1/capacitor_5_2/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.98f
C254 cp2_buffer_5stage_1/cp2_buffer1_1/charge_pump_0/capacitors_5_1/capacitor_5_2/buffer_digital_1/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.58f
C255 cp2_buffer_5stage_1/cp2_buffer1_1/charge_pump_0/capacitors_5_1/capacitor_5_1/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.34f
C256 cp2_buffer_5stage_1/cp2_buffer1_1/charge_pump_0/capacitors_5_1/capacitor_5_1/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.98f
C257 cp2_buffer_5stage_1/cp2_buffer1_1/charge_pump_0/capacitors_5_1/capacitor_5_1/buffer_digital_1/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.58f
C258 cp2_buffer_5stage_1/cp2_buffer1_1/charge_pump_0/capacitors_5_1/capacitor_5_0/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.34f
C259 cp2_buffer_5stage_1/cp2_buffer1_1/charge_pump_0/capacitors_5_1/capacitor_5_0/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.98f
C260 cp2_buffer_5stage_1/cp2_buffer1_1/charge_pump_0/capacitors_5_1/capacitor_5_0/buffer_digital_1/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.58f
C261 cp2_buffer_5stage_1/cp2_buffer1_1/charge_pump_0/input2 cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 14.4f
C262 cp2_buffer_5stage_1/cp2_buffer1_1/charge_pump_0/capacitors_5_1/capacitor_5_7/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.34f
C263 cp2_buffer_5stage_1/cp2_buffer1_1/charge_pump_0/clkb cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 84f
C264 cp2_buffer_5stage_1/cp2_buffer1_1/charge_pump_0/capacitors_5_1/capacitor_5_7/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.98f
C265 cp2_buffer_5stage_1/cp2_buffer1_1/charge_pump_0/capacitors_5_1/capacitor_5_7/buffer_digital_1/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.58f
C266 cp2_buffer_5stage_1/cp2_buffer1_1/charge_pump_0/capacitors_5_1/capacitor_5_6/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.34f
C267 cp2_buffer_5stage_1/cp2_buffer1_1/charge_pump_0/capacitors_5_1/capacitor_5_6/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.98f
C268 cp2_buffer_5stage_1/cp2_buffer1_1/charge_pump_0/capacitors_5_1/capacitor_5_6/buffer_digital_1/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.58f
C269 cp2_buffer_5stage_1/cp2_buffer1_1/charge_pump_0/capacitors_5_1/capacitor_5_5/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.34f
C270 cp2_buffer_5stage_1/cp2_buffer1_1/charge_pump_0/capacitors_5_1/capacitor_5_5/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.98f
C271 cp2_buffer_5stage_1/cp2_buffer1_1/charge_pump_0/capacitors_5_1/capacitor_5_5/buffer_digital_1/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.58f
C272 cp2_buffer_5stage_1/cp2_buffer1_1/charge_pump_0/g1 cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.63f
C273 cp2_buffer_5stage_1/cp2_buffer1_0/charge_pump_0/vs cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 50.2f
C274 cp2_buffer_5stage_1/cp2_buffer1_0/charge_pump_0/clock_0/a_2432_n962# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 8.68f **FLOATING
C275 cp2_buffer_5stage_1/cp2_buffer1_0/charge_pump_0/clock_0/a_2020_n482# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.57f **FLOATING
C276 cp2_buffer_5stage_1/cp2_buffer1_0/charge_pump_0/clock_0/a_344_102# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.81f
C277 cp2_buffer_5stage_1/cp2_buffer1_0/charge_pump_0/clock_0/a_2402_572# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.17f
C278 cp2_buffer_5stage_1/cp2_buffer1_0/charge_pump_0/clock_0/a_344_n986# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.38f
C279 cp2_buffer_5stage_1/cp2_buffer2_0/buffer_digital_2/i cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 7.99f
C280 cp2_buffer_5stage_1/cp2_buffer1_0/charge_pump_0/clock_0/a_3246_118# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 6.83f
C281 cp2_buffer_5stage_1/cp2_buffer1_0/charge_pump_0/g2 cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.44f
C282 cp2_buffer_5stage_1/cp2_buffer1_0/charge_pump_0/capacitors_5_0/capacitor_5_4/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.34f
C283 cp2_buffer_5stage_1/cp2_buffer1_0/charge_pump_0/capacitors_5_0/capacitor_5_4/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.98f
C284 cp2_buffer_5stage_1/cp2_buffer1_0/charge_pump_0/capacitors_5_0/capacitor_5_4/buffer_digital_1/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.58f
C285 cp2_buffer_5stage_1/cp2_buffer1_0/charge_pump_0/capacitors_5_0/capacitor_5_3/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.34f
C286 cp2_buffer_5stage_1/cp2_buffer1_0/charge_pump_0/capacitors_5_0/capacitor_5_3/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.98f
C287 cp2_buffer_5stage_1/cp2_buffer1_0/charge_pump_0/capacitors_5_0/capacitor_5_3/buffer_digital_1/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.58f
C288 scanchain_0/data_out[3] cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 35.7f
C289 cp2_buffer_5stage_1/cp2_buffer1_0/charge_pump_0/capacitors_5_0/capacitor_5_2/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.34f
C290 cp2_buffer_5stage_1/cp2_buffer1_0/charge_pump_0/capacitors_5_0/capacitor_5_2/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.98f
C291 cp2_buffer_5stage_1/cp2_buffer1_0/charge_pump_0/capacitors_5_0/capacitor_5_2/buffer_digital_1/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.58f
C292 cp2_buffer_5stage_1/cp2_buffer1_0/charge_pump_0/capacitors_5_0/capacitor_5_1/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.34f
C293 cp2_buffer_5stage_1/cp2_buffer1_0/charge_pump_0/capacitors_5_0/capacitor_5_1/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.98f
C294 cp2_buffer_5stage_1/cp2_buffer1_0/charge_pump_0/capacitors_5_0/capacitor_5_1/buffer_digital_1/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.58f
C295 cp2_buffer_5stage_1/cp2_buffer1_0/charge_pump_0/capacitors_5_0/capacitor_5_0/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.34f
C296 cp2_buffer_5stage_1/cp2_buffer1_0/charge_pump_0/capacitors_5_0/capacitor_5_0/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.98f
C297 cp2_buffer_5stage_1/cp2_buffer1_0/charge_pump_0/capacitors_5_0/capacitor_5_0/buffer_digital_1/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.58f
C298 cp2_buffer_5stage_1/cp2_buffer1_0/charge_pump_0/input1 cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 15f
C299 cp2_buffer_5stage_1/cp2_buffer1_0/charge_pump_0/capacitors_5_0/capacitor_5_7/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.34f
C300 cp2_buffer_5stage_1/cp2_buffer1_0/charge_pump_0/clk cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 82.2f
C301 scanchain_0/VDD cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 7.91p
C302 cp2_buffer_5stage_1/cp2_buffer1_0/charge_pump_0/capacitors_5_0/capacitor_5_7/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.98f
C303 cp2_buffer_5stage_1/cp2_buffer1_0/charge_pump_0/capacitors_5_0/capacitor_5_7/buffer_digital_1/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.58f
C304 cp2_buffer_5stage_1/cp2_buffer1_0/charge_pump_0/capacitors_5_0/capacitor_5_6/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.34f
C305 cp2_buffer_5stage_1/cp2_buffer1_0/charge_pump_0/capacitors_5_0/capacitor_5_6/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.98f
C306 cp2_buffer_5stage_1/cp2_buffer1_0/charge_pump_0/capacitors_5_0/capacitor_5_6/buffer_digital_1/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.58f
C307 cp2_buffer_5stage_1/cp2_buffer1_0/charge_pump_0/capacitors_5_0/capacitor_5_5/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.34f
C308 cp2_buffer_5stage_1/cp2_buffer1_0/charge_pump_0/capacitors_5_0/capacitor_5_5/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.98f
C309 cp2_buffer_5stage_1/cp2_buffer1_0/charge_pump_0/capacitors_5_0/capacitor_5_5/buffer_digital_1/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.58f
C310 cp2_buffer_5stage_1/cp2_buffer1_0/charge_pump_0/capacitors_5_1/capacitor_5_4/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.34f
C311 cp2_buffer_5stage_1/cp2_buffer1_0/charge_pump_0/capacitors_5_1/capacitor_5_4/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.98f
C312 cp2_buffer_5stage_1/cp2_buffer1_0/charge_pump_0/capacitors_5_1/capacitor_5_4/buffer_digital_1/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.58f
C313 cp2_buffer_5stage_1/cp2_buffer1_0/charge_pump_0/capacitors_5_1/capacitor_5_3/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.34f
C314 cp2_buffer_5stage_1/cp2_buffer1_0/charge_pump_0/capacitors_5_1/capacitor_5_3/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.98f
C315 cp2_buffer_5stage_1/cp2_buffer1_0/charge_pump_0/capacitors_5_1/capacitor_5_3/buffer_digital_1/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.58f
C316 cp2_buffer_5stage_1/cp2_buffer1_0/charge_pump_0/capacitors_5_1/capacitor_5_2/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.34f
C317 cp2_buffer_5stage_1/cp2_buffer1_0/charge_pump_0/capacitors_5_1/capacitor_5_2/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.98f
C318 cp2_buffer_5stage_1/cp2_buffer1_0/charge_pump_0/capacitors_5_1/capacitor_5_2/buffer_digital_1/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.58f
C319 cp2_buffer_5stage_1/cp2_buffer1_0/charge_pump_0/capacitors_5_1/capacitor_5_1/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.34f
C320 cp2_buffer_5stage_1/cp2_buffer1_0/charge_pump_0/capacitors_5_1/capacitor_5_1/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.98f
C321 cp2_buffer_5stage_1/cp2_buffer1_0/charge_pump_0/capacitors_5_1/capacitor_5_1/buffer_digital_1/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.58f
C322 cp2_buffer_5stage_1/cp2_buffer1_0/charge_pump_0/capacitors_5_1/capacitor_5_0/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.34f
C323 cp2_buffer_5stage_1/cp2_buffer1_0/charge_pump_0/capacitors_5_1/capacitor_5_0/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.98f
C324 cp2_buffer_5stage_1/cp2_buffer1_0/charge_pump_0/capacitors_5_1/capacitor_5_0/buffer_digital_1/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.58f
C325 cp2_buffer_5stage_1/cp2_buffer1_0/charge_pump_0/input2 cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 14.4f
C326 cp2_buffer_5stage_1/cp2_buffer1_0/charge_pump_0/capacitors_5_1/capacitor_5_7/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.34f
C327 cp2_buffer_5stage_1/cp2_buffer1_0/charge_pump_0/clkb cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 84f
C328 cp2_buffer_5stage_1/cp2_buffer1_0/charge_pump_0/capacitors_5_1/capacitor_5_7/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.98f
C329 cp2_buffer_5stage_1/cp2_buffer1_0/charge_pump_0/capacitors_5_1/capacitor_5_7/buffer_digital_1/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.58f
C330 cp2_buffer_5stage_1/cp2_buffer1_0/charge_pump_0/capacitors_5_1/capacitor_5_6/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.34f
C331 cp2_buffer_5stage_1/cp2_buffer1_0/charge_pump_0/capacitors_5_1/capacitor_5_6/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.98f
C332 cp2_buffer_5stage_1/cp2_buffer1_0/charge_pump_0/capacitors_5_1/capacitor_5_6/buffer_digital_1/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.58f
C333 cp2_buffer_5stage_1/cp2_buffer1_0/charge_pump_0/capacitors_5_1/capacitor_5_5/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.34f
C334 cp2_buffer_5stage_1/cp2_buffer1_0/charge_pump_0/capacitors_5_1/capacitor_5_5/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.98f
C335 cp2_buffer_5stage_1/cp2_buffer1_0/charge_pump_0/capacitors_5_1/capacitor_5_5/buffer_digital_1/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.58f
C336 cp2_buffer_5stage_1/cp2_buffer1_0/charge_pump_0/g1 cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.63f
C337 cp2_buffer_5stage_0/cp2_buffer1_1/charge_pump_0/vin cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 23f
C338 cp2_buffer_5stage_0/cp2_buffer2_1/charge_pump_reverse_0/clock_0/a_2432_n962# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 8.68f **FLOATING
C339 cp2_buffer_5stage_0/cp2_buffer2_1/charge_pump_reverse_0/clock_0/a_2020_n482# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.57f **FLOATING
C340 cp2_buffer_5stage_0/cp2_buffer2_1/charge_pump_reverse_0/clock_0/a_344_102# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.81f
C341 cp2_buffer_5stage_0/cp2_buffer2_1/charge_pump_reverse_0/clock_0/a_2402_572# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.17f
C342 cp2_buffer_5stage_0/cp2_buffer2_1/charge_pump_reverse_0/clock_0/a_344_n986# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.38f
C343 cp2_buffer_5stage_0/cp2_buffer1_2/buffer_digital_1/i cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 7.37f
C344 cp2_buffer_5stage_0/cp2_buffer2_1/charge_pump_reverse_0/clock_0/a_3246_118# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 6.83f
C345 cp2_buffer_5stage_0/cp2_buffer2_1/charge_pump_reverse_0/nmos_dnw3_0/clkb cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.23f
C346 cp2_buffer_5stage_0/cp2_buffer2_1/charge_pump_reverse_0/capacitors_5_0/capacitor_5_4/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.34f
C347 cp2_buffer_5stage_0/cp2_buffer2_1/charge_pump_reverse_0/capacitors_5_0/capacitor_5_4/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.98f
C348 cp2_buffer_5stage_0/cp2_buffer2_1/charge_pump_reverse_0/capacitors_5_0/capacitor_5_4/buffer_digital_1/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.58f
C349 cp2_buffer_5stage_0/cp2_buffer2_1/charge_pump_reverse_0/capacitors_5_0/capacitor_5_3/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.34f
C350 cp2_buffer_5stage_0/cp2_buffer2_1/charge_pump_reverse_0/capacitors_5_0/capacitor_5_3/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.98f
C351 cp2_buffer_5stage_0/cp2_buffer2_1/charge_pump_reverse_0/capacitors_5_0/capacitor_5_3/buffer_digital_1/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.58f
C352 cp2_buffer_5stage_0/cp2_buffer2_1/charge_pump_reverse_0/capacitors_5_0/capacitor_5_2/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.34f
C353 cp2_buffer_5stage_0/cp2_buffer2_1/charge_pump_reverse_0/capacitors_5_0/capacitor_5_2/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.98f
C354 cp2_buffer_5stage_0/cp2_buffer2_1/charge_pump_reverse_0/capacitors_5_0/capacitor_5_2/buffer_digital_1/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.58f
C355 cp2_buffer_5stage_0/cp2_buffer2_1/charge_pump_reverse_0/capacitors_5_0/capacitor_5_1/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.34f
C356 cp2_buffer_5stage_0/cp2_buffer2_1/charge_pump_reverse_0/capacitors_5_0/capacitor_5_1/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.98f
C357 cp2_buffer_5stage_0/cp2_buffer2_1/charge_pump_reverse_0/capacitors_5_0/capacitor_5_1/buffer_digital_1/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.58f
C358 cp2_buffer_5stage_0/cp2_buffer2_1/charge_pump_reverse_0/capacitors_5_0/capacitor_5_0/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.34f
C359 cp2_buffer_5stage_0/cp2_buffer2_1/charge_pump_reverse_0/capacitors_5_0/capacitor_5_0/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.98f
C360 cp2_buffer_5stage_0/cp2_buffer2_1/charge_pump_reverse_0/capacitors_5_0/capacitor_5_0/buffer_digital_1/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.58f
C361 cp2_buffer_5stage_0/cp2_buffer2_1/charge_pump_reverse_0/nmos_dnw3_0/out1 cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 15.1f
C362 cp2_buffer_5stage_0/cp2_buffer2_1/charge_pump_reverse_0/capacitors_5_0/capacitor_5_7/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.34f
C363 cp2_buffer_5stage_0/cp2_buffer2_1/charge_pump_reverse_0/clock_0/clkb cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 90.9f
C364 cp2_buffer_5stage_0/cp2_buffer2_1/charge_pump_reverse_0/capacitors_5_0/capacitor_5_7/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.98f
C365 cp2_buffer_5stage_0/cp2_buffer2_1/charge_pump_reverse_0/capacitors_5_0/capacitor_5_7/buffer_digital_1/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.58f
C366 cp2_buffer_5stage_0/cp2_buffer2_1/charge_pump_reverse_0/capacitors_5_0/capacitor_5_6/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.34f
C367 cp2_buffer_5stage_0/cp2_buffer2_1/charge_pump_reverse_0/capacitors_5_0/capacitor_5_6/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.98f
C368 cp2_buffer_5stage_0/cp2_buffer2_1/charge_pump_reverse_0/capacitors_5_0/capacitor_5_6/buffer_digital_1/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.58f
C369 cp2_buffer_5stage_0/cp2_buffer2_1/charge_pump_reverse_0/capacitors_5_0/capacitor_5_5/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.34f
C370 cp2_buffer_5stage_0/cp2_buffer2_1/charge_pump_reverse_0/capacitors_5_0/capacitor_5_5/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.98f
C371 cp2_buffer_5stage_0/cp2_buffer2_1/charge_pump_reverse_0/capacitors_5_0/capacitor_5_5/buffer_digital_1/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.58f
C372 cp2_buffer_5stage_0/cp2_buffer2_1/charge_pump_reverse_0/capacitors_5_1/capacitor_5_4/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.34f
C373 cp2_buffer_5stage_0/cp2_buffer2_1/charge_pump_reverse_0/capacitors_5_1/capacitor_5_4/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.98f
C374 cp2_buffer_5stage_0/cp2_buffer2_1/charge_pump_reverse_0/capacitors_5_1/capacitor_5_4/buffer_digital_1/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.58f
C375 cp2_buffer_5stage_0/cp2_buffer2_1/charge_pump_reverse_0/capacitors_5_1/capacitor_5_3/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.34f
C376 cp2_buffer_5stage_0/cp2_buffer2_1/charge_pump_reverse_0/capacitors_5_1/capacitor_5_3/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.98f
C377 cp2_buffer_5stage_0/cp2_buffer2_1/charge_pump_reverse_0/capacitors_5_1/capacitor_5_3/buffer_digital_1/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.58f
C378 cp2_buffer_5stage_0/cp2_buffer2_1/charge_pump_reverse_0/capacitors_5_1/capacitor_5_2/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.34f
C379 cp2_buffer_5stage_0/cp2_buffer2_1/charge_pump_reverse_0/capacitors_5_1/capacitor_5_2/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.98f
C380 cp2_buffer_5stage_0/cp2_buffer2_1/charge_pump_reverse_0/capacitors_5_1/capacitor_5_2/buffer_digital_1/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.58f
C381 cp2_buffer_5stage_0/cp2_buffer2_1/charge_pump_reverse_0/capacitors_5_1/capacitor_5_1/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.34f
C382 cp2_buffer_5stage_0/cp2_buffer2_1/charge_pump_reverse_0/capacitors_5_1/capacitor_5_1/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.98f
C383 cp2_buffer_5stage_0/cp2_buffer2_1/charge_pump_reverse_0/capacitors_5_1/capacitor_5_1/buffer_digital_1/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.58f
C384 cp2_buffer_5stage_0/cp2_buffer2_1/charge_pump_reverse_0/capacitors_5_1/capacitor_5_0/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.34f
C385 cp2_buffer_5stage_0/cp2_buffer2_1/charge_pump_reverse_0/capacitors_5_1/capacitor_5_0/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.98f
C386 cp2_buffer_5stage_0/cp2_buffer2_1/charge_pump_reverse_0/capacitors_5_1/capacitor_5_0/buffer_digital_1/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.58f
C387 cp2_buffer_5stage_0/cp2_buffer2_1/charge_pump_reverse_0/nmos_dnw3_0/out2 cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 14.8f
C388 cp2_buffer_5stage_0/cp2_buffer2_1/charge_pump_reverse_0/capacitors_5_1/capacitor_5_7/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.34f
C389 cp2_buffer_5stage_0/cp2_buffer2_1/charge_pump_reverse_0/clock_0/clk cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 84.5f
C390 cp2_buffer_5stage_0/cp2_buffer2_1/charge_pump_reverse_0/capacitors_5_1/capacitor_5_7/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.98f
C391 cp2_buffer_5stage_0/cp2_buffer2_1/charge_pump_reverse_0/capacitors_5_1/capacitor_5_7/buffer_digital_1/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.58f
C392 cp2_buffer_5stage_0/cp2_buffer2_1/charge_pump_reverse_0/capacitors_5_1/capacitor_5_6/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.34f
C393 cp2_buffer_5stage_0/cp2_buffer2_1/charge_pump_reverse_0/capacitors_5_1/capacitor_5_6/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.98f
C394 cp2_buffer_5stage_0/cp2_buffer2_1/charge_pump_reverse_0/capacitors_5_1/capacitor_5_6/buffer_digital_1/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.58f
C395 cp2_buffer_5stage_0/cp2_buffer2_1/charge_pump_reverse_0/capacitors_5_1/capacitor_5_5/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.34f
C396 cp2_buffer_5stage_0/cp2_buffer2_1/charge_pump_reverse_0/capacitors_5_1/capacitor_5_5/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.98f
C397 cp2_buffer_5stage_0/cp2_buffer2_1/charge_pump_reverse_0/capacitors_5_1/capacitor_5_5/buffer_digital_1/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.58f
C398 cp2_buffer_5stage_0/cp2_buffer2_1/charge_pump_reverse_0/nmos_dnw3_0/clk cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.43f
C399 cp2_buffer_5stage_0/cp2_buffer1_0/charge_pump_0/vin cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 33.4f
C400 cp2_buffer_5stage_0/cp2_buffer2_0/charge_pump_reverse_0/clock_0/a_2432_n962# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 8.68f **FLOATING
C401 cp2_buffer_5stage_0/cp2_buffer2_0/charge_pump_reverse_0/clock_0/a_2020_n482# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.57f **FLOATING
C402 cp2_buffer_5stage_0/cp2_buffer2_0/charge_pump_reverse_0/clock_0/a_344_102# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.81f
C403 cp2_buffer_5stage_0/cp2_buffer2_0/charge_pump_reverse_0/clock_0/a_2402_572# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.17f
C404 cp2_buffer_5stage_0/cp2_buffer2_0/charge_pump_reverse_0/clock_0/a_344_n986# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.38f
C405 cp2_buffer_5stage_0/cp2_buffer1_1/buffer_digital_1/i cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 7.27f
C406 cp2_buffer_5stage_0/cp2_buffer2_0/charge_pump_reverse_0/clock_0/a_3246_118# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 6.83f
C407 cp2_buffer_5stage_0/cp2_buffer2_0/charge_pump_reverse_0/nmos_dnw3_0/clkb cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.23f
C408 cp2_buffer_5stage_0/cp2_buffer2_0/charge_pump_reverse_0/capacitors_5_0/capacitor_5_4/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.34f
C409 cp2_buffer_5stage_0/cp2_buffer2_0/charge_pump_reverse_0/capacitors_5_0/capacitor_5_4/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.98f
C410 cp2_buffer_5stage_0/cp2_buffer2_0/charge_pump_reverse_0/capacitors_5_0/capacitor_5_4/buffer_digital_1/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.58f
C411 cp2_buffer_5stage_0/cp2_buffer2_0/charge_pump_reverse_0/capacitors_5_0/capacitor_5_3/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.34f
C412 cp2_buffer_5stage_0/cp2_buffer2_0/charge_pump_reverse_0/capacitors_5_0/capacitor_5_3/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.98f
C413 cp2_buffer_5stage_0/cp2_buffer2_0/charge_pump_reverse_0/capacitors_5_0/capacitor_5_3/buffer_digital_1/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.58f
C414 cp2_buffer_5stage_0/cp2_buffer2_0/charge_pump_reverse_0/capacitors_5_0/capacitor_5_2/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.34f
C415 cp2_buffer_5stage_0/cp2_buffer2_0/charge_pump_reverse_0/capacitors_5_0/capacitor_5_2/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.98f
C416 cp2_buffer_5stage_0/cp2_buffer2_0/charge_pump_reverse_0/capacitors_5_0/capacitor_5_2/buffer_digital_1/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.58f
C417 cp2_buffer_5stage_0/cp2_buffer2_0/charge_pump_reverse_0/capacitors_5_0/capacitor_5_1/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.34f
C418 cp2_buffer_5stage_0/cp2_buffer2_0/charge_pump_reverse_0/capacitors_5_0/capacitor_5_1/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.98f
C419 cp2_buffer_5stage_0/cp2_buffer2_0/charge_pump_reverse_0/capacitors_5_0/capacitor_5_1/buffer_digital_1/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.58f
C420 cp2_buffer_5stage_0/cp2_buffer2_0/charge_pump_reverse_0/capacitors_5_0/capacitor_5_0/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.34f
C421 cp2_buffer_5stage_0/cp2_buffer2_0/charge_pump_reverse_0/capacitors_5_0/capacitor_5_0/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.98f
C422 cp2_buffer_5stage_0/cp2_buffer2_0/charge_pump_reverse_0/capacitors_5_0/capacitor_5_0/buffer_digital_1/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.58f
C423 cp2_buffer_5stage_0/cp2_buffer2_0/charge_pump_reverse_0/nmos_dnw3_0/out1 cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 15.1f
C424 cp2_buffer_5stage_0/cp2_buffer2_0/charge_pump_reverse_0/capacitors_5_0/capacitor_5_7/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.34f
C425 cp2_buffer_5stage_0/cp2_buffer2_0/charge_pump_reverse_0/clock_0/clkb cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 90.9f
C426 cp2_buffer_5stage_0/cp2_buffer2_0/charge_pump_reverse_0/capacitors_5_0/capacitor_5_7/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.98f
C427 cp2_buffer_5stage_0/cp2_buffer2_0/charge_pump_reverse_0/capacitors_5_0/capacitor_5_7/buffer_digital_1/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.58f
C428 cp2_buffer_5stage_0/cp2_buffer2_0/charge_pump_reverse_0/capacitors_5_0/capacitor_5_6/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.34f
C429 cp2_buffer_5stage_0/cp2_buffer2_0/charge_pump_reverse_0/capacitors_5_0/capacitor_5_6/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.98f
C430 cp2_buffer_5stage_0/cp2_buffer2_0/charge_pump_reverse_0/capacitors_5_0/capacitor_5_6/buffer_digital_1/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.58f
C431 cp2_buffer_5stage_0/cp2_buffer2_0/charge_pump_reverse_0/capacitors_5_0/capacitor_5_5/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.34f
C432 cp2_buffer_5stage_0/cp2_buffer2_0/charge_pump_reverse_0/capacitors_5_0/capacitor_5_5/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.98f
C433 cp2_buffer_5stage_0/cp2_buffer2_0/charge_pump_reverse_0/capacitors_5_0/capacitor_5_5/buffer_digital_1/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.58f
C434 cp2_buffer_5stage_0/cp2_buffer2_0/charge_pump_reverse_0/capacitors_5_1/capacitor_5_4/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.34f
C435 cp2_buffer_5stage_0/cp2_buffer2_0/charge_pump_reverse_0/capacitors_5_1/capacitor_5_4/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.98f
C436 cp2_buffer_5stage_0/cp2_buffer2_0/charge_pump_reverse_0/capacitors_5_1/capacitor_5_4/buffer_digital_1/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.58f
C437 cp2_buffer_5stage_0/cp2_buffer2_0/charge_pump_reverse_0/capacitors_5_1/capacitor_5_3/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.34f
C438 cp2_buffer_5stage_0/cp2_buffer2_0/charge_pump_reverse_0/capacitors_5_1/capacitor_5_3/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.98f
C439 cp2_buffer_5stage_0/cp2_buffer2_0/charge_pump_reverse_0/capacitors_5_1/capacitor_5_3/buffer_digital_1/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.58f
C440 cp2_buffer_5stage_0/cp2_buffer2_0/charge_pump_reverse_0/capacitors_5_1/capacitor_5_2/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.34f
C441 cp2_buffer_5stage_0/cp2_buffer2_0/charge_pump_reverse_0/capacitors_5_1/capacitor_5_2/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.98f
C442 cp2_buffer_5stage_0/cp2_buffer2_0/charge_pump_reverse_0/capacitors_5_1/capacitor_5_2/buffer_digital_1/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.58f
C443 cp2_buffer_5stage_0/cp2_buffer2_0/charge_pump_reverse_0/capacitors_5_1/capacitor_5_1/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.34f
C444 cp2_buffer_5stage_0/cp2_buffer2_0/charge_pump_reverse_0/capacitors_5_1/capacitor_5_1/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.98f
C445 cp2_buffer_5stage_0/cp2_buffer2_0/charge_pump_reverse_0/capacitors_5_1/capacitor_5_1/buffer_digital_1/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.58f
C446 cp2_buffer_5stage_0/cp2_buffer2_0/charge_pump_reverse_0/capacitors_5_1/capacitor_5_0/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.34f
C447 cp2_buffer_5stage_0/cp2_buffer2_0/charge_pump_reverse_0/capacitors_5_1/capacitor_5_0/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.98f
C448 cp2_buffer_5stage_0/cp2_buffer2_0/charge_pump_reverse_0/capacitors_5_1/capacitor_5_0/buffer_digital_1/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.58f
C449 scanchain_0/data_out[0] cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 52.6f
C450 cp2_buffer_5stage_0/cp2_buffer2_0/charge_pump_reverse_0/nmos_dnw3_0/out2 cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 14.8f
C451 cp2_buffer_5stage_0/cp2_buffer2_0/charge_pump_reverse_0/capacitors_5_1/capacitor_5_7/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.34f
C452 cp2_buffer_5stage_0/cp2_buffer2_0/charge_pump_reverse_0/clock_0/clk cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 84.5f
C453 cp2_buffer_5stage_0/cp2_buffer2_0/charge_pump_reverse_0/capacitors_5_1/capacitor_5_7/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.98f
C454 cp2_buffer_5stage_0/cp2_buffer2_0/charge_pump_reverse_0/capacitors_5_1/capacitor_5_7/buffer_digital_1/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.58f
C455 cp2_buffer_5stage_0/cp2_buffer2_0/charge_pump_reverse_0/capacitors_5_1/capacitor_5_6/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.34f
C456 cp2_buffer_5stage_0/cp2_buffer2_0/charge_pump_reverse_0/capacitors_5_1/capacitor_5_6/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.98f
C457 cp2_buffer_5stage_0/cp2_buffer2_0/charge_pump_reverse_0/capacitors_5_1/capacitor_5_6/buffer_digital_1/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.58f
C458 cp2_buffer_5stage_0/cp2_buffer2_0/charge_pump_reverse_0/capacitors_5_1/capacitor_5_5/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.34f
C459 cp2_buffer_5stage_0/cp2_buffer2_0/charge_pump_reverse_0/capacitors_5_1/capacitor_5_5/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.98f
C460 cp2_buffer_5stage_0/cp2_buffer2_0/charge_pump_reverse_0/capacitors_5_1/capacitor_5_5/buffer_digital_1/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.58f
C461 cp2_buffer_5stage_0/cp2_buffer2_0/charge_pump_reverse_0/nmos_dnw3_0/clk cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.43f
C462 cp2_buffer_5stage_0/cp2_buffer1_2/charge_pump_0/vin cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 3.29f
C463 cp2_buffer_5stage_0/cp2_buffer1_2/charge_pump_0/clock_0/a_2432_n962# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 8.68f **FLOATING
C464 cp2_buffer_5stage_0/cp2_buffer1_2/charge_pump_0/clock_0/a_2020_n482# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.57f **FLOATING
C465 cp2_buffer_5stage_0/cp2_buffer1_2/charge_pump_0/clock_0/a_344_102# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.81f
C466 cp2_buffer_5stage_0/cp2_buffer1_2/charge_pump_0/clock_0/a_2402_572# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.17f
C467 cp2_buffer_5stage_0/cp2_buffer1_2/charge_pump_0/clock_0/a_344_n986# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.38f
C468 cp2_buffer_5stage_0/cp2_buffer1_2/buffer_digital_0/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.95f
C469 cp2_buffer_5stage_0/cp2_buffer1_2/charge_pump_0/clock_0/a_3246_118# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 6.83f
C470 cp2_buffer_5stage_0/cp2_buffer1_2/charge_pump_0/g2 cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.44f
C471 cp2_buffer_5stage_0/cp2_buffer1_2/charge_pump_0/capacitors_5_0/capacitor_5_4/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.34f
C472 cp2_buffer_5stage_0/cp2_buffer1_2/charge_pump_0/capacitors_5_0/capacitor_5_4/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.98f
C473 cp2_buffer_5stage_0/cp2_buffer1_2/charge_pump_0/capacitors_5_0/capacitor_5_4/buffer_digital_1/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.58f
C474 cp2_buffer_5stage_0/cp2_buffer1_2/charge_pump_0/capacitors_5_0/capacitor_5_3/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.34f
C475 cp2_buffer_5stage_0/cp2_buffer1_2/charge_pump_0/capacitors_5_0/capacitor_5_3/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.98f
C476 cp2_buffer_5stage_0/cp2_buffer1_2/charge_pump_0/capacitors_5_0/capacitor_5_3/buffer_digital_1/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.58f
C477 cp2_buffer_5stage_0/cp2_buffer1_2/charge_pump_0/capacitors_5_0/capacitor_5_2/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.34f
C478 cp2_buffer_5stage_0/cp2_buffer1_2/charge_pump_0/capacitors_5_0/capacitor_5_2/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.98f
C479 cp2_buffer_5stage_0/cp2_buffer1_2/charge_pump_0/capacitors_5_0/capacitor_5_2/buffer_digital_1/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.58f
C480 cp2_buffer_5stage_0/cp2_buffer1_2/charge_pump_0/capacitors_5_0/capacitor_5_1/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.34f
C481 cp2_buffer_5stage_0/cp2_buffer1_2/charge_pump_0/capacitors_5_0/capacitor_5_1/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.98f
C482 cp2_buffer_5stage_0/cp2_buffer1_2/charge_pump_0/capacitors_5_0/capacitor_5_1/buffer_digital_1/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.58f
C483 cp2_buffer_5stage_0/cp2_buffer1_2/charge_pump_0/capacitors_5_0/capacitor_5_0/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.34f
C484 cp2_buffer_5stage_0/cp2_buffer1_2/charge_pump_0/capacitors_5_0/capacitor_5_0/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.98f
C485 cp2_buffer_5stage_0/cp2_buffer1_2/charge_pump_0/capacitors_5_0/capacitor_5_0/buffer_digital_1/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.58f
C486 cp2_buffer_5stage_0/cp2_buffer1_2/charge_pump_0/input1 cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 15f
C487 cp2_buffer_5stage_0/cp2_buffer1_2/charge_pump_0/capacitors_5_0/capacitor_5_7/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.34f
C488 cp2_buffer_5stage_0/cp2_buffer1_2/charge_pump_0/clk cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 82.3f
C489 cp2_buffer_5stage_0/cp2_buffer1_2/charge_pump_0/capacitors_5_0/capacitor_5_7/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.98f
C490 cp2_buffer_5stage_0/cp2_buffer1_2/charge_pump_0/capacitors_5_0/capacitor_5_7/buffer_digital_1/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.58f
C491 cp2_buffer_5stage_0/cp2_buffer1_2/charge_pump_0/capacitors_5_0/capacitor_5_6/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.34f
C492 cp2_buffer_5stage_0/cp2_buffer1_2/charge_pump_0/capacitors_5_0/capacitor_5_6/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.98f
C493 cp2_buffer_5stage_0/cp2_buffer1_2/charge_pump_0/capacitors_5_0/capacitor_5_6/buffer_digital_1/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.58f
C494 cp2_buffer_5stage_0/cp2_buffer1_2/charge_pump_0/capacitors_5_0/capacitor_5_5/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.34f
C495 cp2_buffer_5stage_0/cp2_buffer1_2/charge_pump_0/capacitors_5_0/capacitor_5_5/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.98f
C496 cp2_buffer_5stage_0/cp2_buffer1_2/charge_pump_0/capacitors_5_0/capacitor_5_5/buffer_digital_1/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.58f
C497 cp2_buffer_5stage_0/cp2_buffer1_2/charge_pump_0/capacitors_5_1/capacitor_5_4/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.34f
C498 cp2_buffer_5stage_0/cp2_buffer1_2/charge_pump_0/capacitors_5_1/capacitor_5_4/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.98f
C499 cp2_buffer_5stage_0/cp2_buffer1_2/charge_pump_0/capacitors_5_1/capacitor_5_4/buffer_digital_1/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.58f
C500 cp2_buffer_5stage_0/cp2_buffer1_2/charge_pump_0/capacitors_5_1/capacitor_5_3/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.34f
C501 cp2_buffer_5stage_0/cp2_buffer1_2/charge_pump_0/capacitors_5_1/capacitor_5_3/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.98f
C502 cp2_buffer_5stage_0/cp2_buffer1_2/charge_pump_0/capacitors_5_1/capacitor_5_3/buffer_digital_1/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.58f
C503 cp2_buffer_5stage_0/cp2_buffer1_2/charge_pump_0/capacitors_5_1/capacitor_5_2/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.34f
C504 cp2_buffer_5stage_0/cp2_buffer1_2/charge_pump_0/capacitors_5_1/capacitor_5_2/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.98f
C505 cp2_buffer_5stage_0/cp2_buffer1_2/charge_pump_0/capacitors_5_1/capacitor_5_2/buffer_digital_1/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.58f
C506 cp2_buffer_5stage_0/cp2_buffer1_2/charge_pump_0/capacitors_5_1/capacitor_5_1/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.34f
C507 cp2_buffer_5stage_0/cp2_buffer1_2/charge_pump_0/capacitors_5_1/capacitor_5_1/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.98f
C508 cp2_buffer_5stage_0/cp2_buffer1_2/charge_pump_0/capacitors_5_1/capacitor_5_1/buffer_digital_1/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.58f
C509 cp2_buffer_5stage_0/cp2_buffer1_2/charge_pump_0/capacitors_5_1/capacitor_5_0/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.34f
C510 cp2_buffer_5stage_0/cp2_buffer1_2/charge_pump_0/capacitors_5_1/capacitor_5_0/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.98f
C511 cp2_buffer_5stage_0/cp2_buffer1_2/charge_pump_0/capacitors_5_1/capacitor_5_0/buffer_digital_1/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.58f
C512 cp2_buffer_5stage_0/cp2_buffer1_2/charge_pump_0/input2 cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 14.4f
C513 cp2_buffer_5stage_0/cp2_buffer1_2/charge_pump_0/capacitors_5_1/capacitor_5_7/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.34f
C514 cp2_buffer_5stage_0/cp2_buffer1_2/charge_pump_0/clkb cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 84f
C515 cp2_buffer_5stage_0/cp2_buffer1_2/charge_pump_0/capacitors_5_1/capacitor_5_7/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.98f
C516 cp2_buffer_5stage_0/cp2_buffer1_2/charge_pump_0/capacitors_5_1/capacitor_5_7/buffer_digital_1/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.58f
C517 cp2_buffer_5stage_0/cp2_buffer1_2/charge_pump_0/capacitors_5_1/capacitor_5_6/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.34f
C518 cp2_buffer_5stage_0/cp2_buffer1_2/charge_pump_0/capacitors_5_1/capacitor_5_6/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.98f
C519 cp2_buffer_5stage_0/cp2_buffer1_2/charge_pump_0/capacitors_5_1/capacitor_5_6/buffer_digital_1/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.58f
C520 cp2_buffer_5stage_0/cp2_buffer1_2/charge_pump_0/capacitors_5_1/capacitor_5_5/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.34f
C521 cp2_buffer_5stage_0/cp2_buffer1_2/charge_pump_0/capacitors_5_1/capacitor_5_5/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.98f
C522 cp2_buffer_5stage_0/cp2_buffer1_2/charge_pump_0/capacitors_5_1/capacitor_5_5/buffer_digital_1/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.58f
C523 cp2_buffer_5stage_0/cp2_buffer1_2/charge_pump_0/g1 cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.63f
C524 cp2_buffer_5stage_0/cp2_buffer1_1/charge_pump_0/vs cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 24f
C525 cp2_buffer_5stage_0/cp2_buffer1_1/charge_pump_0/clock_0/a_2432_n962# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 8.68f **FLOATING
C526 cp2_buffer_5stage_0/cp2_buffer1_1/charge_pump_0/clock_0/a_2020_n482# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.57f **FLOATING
C527 cp2_buffer_5stage_0/cp2_buffer1_1/charge_pump_0/clock_0/a_344_102# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.81f
C528 cp2_buffer_5stage_0/cp2_buffer1_1/charge_pump_0/clock_0/a_2402_572# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.17f
C529 cp2_buffer_5stage_0/cp2_buffer1_1/charge_pump_0/clock_0/a_344_n986# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.38f
C530 cp2_buffer_5stage_0/cp2_buffer2_1/buffer_digital_2/i cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 6.84f
C531 cp2_buffer_5stage_0/cp2_buffer1_1/charge_pump_0/clock_0/a_3246_118# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 6.83f
C532 cp2_buffer_5stage_0/cp2_buffer1_1/charge_pump_0/g2 cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.44f
C533 cp2_buffer_5stage_0/cp2_buffer1_1/charge_pump_0/capacitors_5_0/capacitor_5_4/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.34f
C534 cp2_buffer_5stage_0/cp2_buffer1_1/charge_pump_0/capacitors_5_0/capacitor_5_4/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.98f
C535 cp2_buffer_5stage_0/cp2_buffer1_1/charge_pump_0/capacitors_5_0/capacitor_5_4/buffer_digital_1/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.58f
C536 cp2_buffer_5stage_0/cp2_buffer1_1/charge_pump_0/capacitors_5_0/capacitor_5_3/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.34f
C537 cp2_buffer_5stage_0/cp2_buffer1_1/charge_pump_0/capacitors_5_0/capacitor_5_3/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.98f
C538 cp2_buffer_5stage_0/cp2_buffer1_1/charge_pump_0/capacitors_5_0/capacitor_5_3/buffer_digital_1/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.58f
C539 cp2_buffer_5stage_0/cp2_buffer1_1/charge_pump_0/capacitors_5_0/capacitor_5_2/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.34f
C540 cp2_buffer_5stage_0/cp2_buffer1_1/charge_pump_0/capacitors_5_0/capacitor_5_2/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.98f
C541 cp2_buffer_5stage_0/cp2_buffer1_1/charge_pump_0/capacitors_5_0/capacitor_5_2/buffer_digital_1/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.58f
C542 cp2_buffer_5stage_0/cp2_buffer1_1/charge_pump_0/capacitors_5_0/capacitor_5_1/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.34f
C543 cp2_buffer_5stage_0/cp2_buffer1_1/charge_pump_0/capacitors_5_0/capacitor_5_1/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.98f
C544 cp2_buffer_5stage_0/cp2_buffer1_1/charge_pump_0/capacitors_5_0/capacitor_5_1/buffer_digital_1/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.58f
C545 scanchain_0/data_out[6] cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 51.9f
C546 cp2_buffer_5stage_0/cp2_buffer1_1/charge_pump_0/capacitors_5_0/capacitor_5_0/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.34f
C547 cp2_buffer_5stage_0/cp2_buffer1_1/charge_pump_0/capacitors_5_0/capacitor_5_0/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.98f
C548 cp2_buffer_5stage_0/cp2_buffer1_1/charge_pump_0/capacitors_5_0/capacitor_5_0/buffer_digital_1/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.58f
C549 cp2_buffer_5stage_0/cp2_buffer1_1/charge_pump_0/input1 cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 15f
C550 cp2_buffer_5stage_0/cp2_buffer1_1/charge_pump_0/capacitors_5_0/capacitor_5_7/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.34f
C551 cp2_buffer_5stage_0/cp2_buffer1_1/charge_pump_0/clk cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 82.3f
C552 cp2_buffer_5stage_0/cp2_buffer1_1/charge_pump_0/capacitors_5_0/capacitor_5_7/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.98f
C553 cp2_buffer_5stage_0/cp2_buffer1_1/charge_pump_0/capacitors_5_0/capacitor_5_7/buffer_digital_1/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.58f
C554 cp2_buffer_5stage_0/cp2_buffer1_1/charge_pump_0/capacitors_5_0/capacitor_5_6/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.34f
C555 cp2_buffer_5stage_0/cp2_buffer1_1/charge_pump_0/capacitors_5_0/capacitor_5_6/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.98f
C556 cp2_buffer_5stage_0/cp2_buffer1_1/charge_pump_0/capacitors_5_0/capacitor_5_6/buffer_digital_1/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.58f
C557 cp2_buffer_5stage_0/cp2_buffer1_1/charge_pump_0/capacitors_5_0/capacitor_5_5/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.34f
C558 cp2_buffer_5stage_0/cp2_buffer1_1/charge_pump_0/capacitors_5_0/capacitor_5_5/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.98f
C559 cp2_buffer_5stage_0/cp2_buffer1_1/charge_pump_0/capacitors_5_0/capacitor_5_5/buffer_digital_1/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.58f
C560 cp2_buffer_5stage_0/cp2_buffer1_1/charge_pump_0/capacitors_5_1/capacitor_5_4/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.34f
C561 cp2_buffer_5stage_0/cp2_buffer1_1/charge_pump_0/capacitors_5_1/capacitor_5_4/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.98f
C562 cp2_buffer_5stage_0/cp2_buffer1_1/charge_pump_0/capacitors_5_1/capacitor_5_4/buffer_digital_1/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.58f
C563 cp2_buffer_5stage_0/cp2_buffer1_1/charge_pump_0/capacitors_5_1/capacitor_5_3/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.34f
C564 cp2_buffer_5stage_0/cp2_buffer1_1/charge_pump_0/capacitors_5_1/capacitor_5_3/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.98f
C565 cp2_buffer_5stage_0/cp2_buffer1_1/charge_pump_0/capacitors_5_1/capacitor_5_3/buffer_digital_1/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.58f
C566 cp2_buffer_5stage_0/cp2_buffer1_1/charge_pump_0/capacitors_5_1/capacitor_5_2/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.34f
C567 cp2_buffer_5stage_0/cp2_buffer1_1/charge_pump_0/capacitors_5_1/capacitor_5_2/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.98f
C568 cp2_buffer_5stage_0/cp2_buffer1_1/charge_pump_0/capacitors_5_1/capacitor_5_2/buffer_digital_1/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.58f
C569 cp2_buffer_5stage_0/cp2_buffer1_1/charge_pump_0/capacitors_5_1/capacitor_5_1/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.34f
C570 cp2_buffer_5stage_0/cp2_buffer1_1/charge_pump_0/capacitors_5_1/capacitor_5_1/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.98f
C571 cp2_buffer_5stage_0/cp2_buffer1_1/charge_pump_0/capacitors_5_1/capacitor_5_1/buffer_digital_1/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.58f
C572 cp2_buffer_5stage_0/cp2_buffer1_1/charge_pump_0/capacitors_5_1/capacitor_5_0/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.34f
C573 cp2_buffer_5stage_0/cp2_buffer1_1/charge_pump_0/capacitors_5_1/capacitor_5_0/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.98f
C574 cp2_buffer_5stage_0/cp2_buffer1_1/charge_pump_0/capacitors_5_1/capacitor_5_0/buffer_digital_1/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.58f
C575 cp2_buffer_5stage_0/cp2_buffer1_1/charge_pump_0/input2 cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 14.4f
C576 cp2_buffer_5stage_0/cp2_buffer1_1/charge_pump_0/capacitors_5_1/capacitor_5_7/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.34f
C577 cp2_buffer_5stage_0/cp2_buffer1_1/charge_pump_0/clkb cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 84f
C578 cp2_buffer_5stage_0/cp2_buffer1_1/charge_pump_0/capacitors_5_1/capacitor_5_7/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.98f
C579 cp2_buffer_5stage_0/cp2_buffer1_1/charge_pump_0/capacitors_5_1/capacitor_5_7/buffer_digital_1/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.58f
C580 cp2_buffer_5stage_0/cp2_buffer1_1/charge_pump_0/capacitors_5_1/capacitor_5_6/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.34f
C581 cp2_buffer_5stage_0/cp2_buffer1_1/charge_pump_0/capacitors_5_1/capacitor_5_6/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.98f
C582 cp2_buffer_5stage_0/cp2_buffer1_1/charge_pump_0/capacitors_5_1/capacitor_5_6/buffer_digital_1/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.58f
C583 cp2_buffer_5stage_0/cp2_buffer1_1/charge_pump_0/capacitors_5_1/capacitor_5_5/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.34f
C584 cp2_buffer_5stage_0/cp2_buffer1_1/charge_pump_0/capacitors_5_1/capacitor_5_5/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.98f
C585 cp2_buffer_5stage_0/cp2_buffer1_1/charge_pump_0/capacitors_5_1/capacitor_5_5/buffer_digital_1/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.58f
C586 cp2_buffer_5stage_0/cp2_buffer1_1/charge_pump_0/g1 cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.63f
C587 cp2_buffer_5stage_0/cp2_buffer1_0/charge_pump_0/clock_0/a_2432_n962# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 8.68f **FLOATING
C588 cp2_buffer_5stage_0/cp2_buffer1_0/charge_pump_0/clock_0/a_2020_n482# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.57f **FLOATING
C589 cp2_buffer_5stage_0/cp2_buffer1_0/charge_pump_0/clock_0/a_344_102# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.81f
C590 cp2_buffer_5stage_0/cp2_buffer1_0/charge_pump_0/clock_0/a_2402_572# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.17f
C591 cp2_buffer_5stage_0/cp2_buffer1_0/charge_pump_0/clock_0/a_344_n986# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.38f
C592 cp2_buffer_5stage_0/cp2_buffer2_0/buffer_digital_2/i cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 7.99f
C593 cp2_buffer_5stage_0/cp2_buffer1_0/charge_pump_0/clock_0/a_3246_118# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 6.83f
C594 cp2_buffer_5stage_0/cp2_buffer1_0/charge_pump_0/g2 cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.44f
C595 cp2_buffer_5stage_0/cp2_buffer1_0/charge_pump_0/capacitors_5_0/capacitor_5_4/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.34f
C596 cp2_buffer_5stage_0/cp2_buffer1_0/charge_pump_0/capacitors_5_0/capacitor_5_4/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.98f
C597 cp2_buffer_5stage_0/cp2_buffer1_0/charge_pump_0/capacitors_5_0/capacitor_5_4/buffer_digital_1/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.58f
C598 cp2_buffer_5stage_0/cp2_buffer1_0/charge_pump_0/capacitors_5_0/capacitor_5_3/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.34f
C599 cp2_buffer_5stage_0/cp2_buffer1_0/charge_pump_0/capacitors_5_0/capacitor_5_3/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.98f
C600 cp2_buffer_5stage_0/cp2_buffer1_0/charge_pump_0/capacitors_5_0/capacitor_5_3/buffer_digital_1/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.58f
C601 scanchain_0/data_out[4] cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 36.9f
C602 cp2_buffer_5stage_0/cp2_buffer1_0/charge_pump_0/capacitors_5_0/capacitor_5_2/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.34f
C603 cp2_buffer_5stage_0/cp2_buffer1_0/charge_pump_0/capacitors_5_0/capacitor_5_2/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.98f
C604 cp2_buffer_5stage_0/cp2_buffer1_0/charge_pump_0/capacitors_5_0/capacitor_5_2/buffer_digital_1/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.58f
C605 cp2_buffer_5stage_0/cp2_buffer1_0/charge_pump_0/capacitors_5_0/capacitor_5_1/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.34f
C606 cp2_buffer_5stage_0/cp2_buffer1_0/charge_pump_0/capacitors_5_0/capacitor_5_1/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.98f
C607 cp2_buffer_5stage_0/cp2_buffer1_0/charge_pump_0/capacitors_5_0/capacitor_5_1/buffer_digital_1/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.58f
C608 cp2_buffer_5stage_0/cp2_buffer1_0/charge_pump_0/capacitors_5_0/capacitor_5_0/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.34f
C609 cp2_buffer_5stage_0/cp2_buffer1_0/charge_pump_0/capacitors_5_0/capacitor_5_0/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.98f
C610 cp2_buffer_5stage_0/cp2_buffer1_0/charge_pump_0/capacitors_5_0/capacitor_5_0/buffer_digital_1/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.58f
C611 cp2_buffer_5stage_0/cp2_buffer1_0/charge_pump_0/input1 cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 15f
C612 cp2_buffer_5stage_0/cp2_buffer1_0/charge_pump_0/capacitors_5_0/capacitor_5_7/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.34f
C613 cp2_buffer_5stage_0/cp2_buffer1_0/charge_pump_0/clk cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 82.3f
C614 cp2_buffer_5stage_0/cp2_buffer1_0/charge_pump_0/capacitors_5_0/capacitor_5_7/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.98f
C615 cp2_buffer_5stage_0/cp2_buffer1_0/charge_pump_0/capacitors_5_0/capacitor_5_7/buffer_digital_1/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.58f
C616 cp2_buffer_5stage_0/cp2_buffer1_0/charge_pump_0/capacitors_5_0/capacitor_5_6/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.34f
C617 cp2_buffer_5stage_0/cp2_buffer1_0/charge_pump_0/capacitors_5_0/capacitor_5_6/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.98f
C618 cp2_buffer_5stage_0/cp2_buffer1_0/charge_pump_0/capacitors_5_0/capacitor_5_6/buffer_digital_1/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.58f
C619 cp2_buffer_5stage_0/cp2_buffer1_0/charge_pump_0/capacitors_5_0/capacitor_5_5/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.34f
C620 cp2_buffer_5stage_0/cp2_buffer1_0/charge_pump_0/capacitors_5_0/capacitor_5_5/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.98f
C621 cp2_buffer_5stage_0/cp2_buffer1_0/charge_pump_0/capacitors_5_0/capacitor_5_5/buffer_digital_1/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.58f
C622 cp2_buffer_5stage_0/cp2_buffer1_0/charge_pump_0/capacitors_5_1/capacitor_5_4/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.34f
C623 cp2_buffer_5stage_0/cp2_buffer1_0/charge_pump_0/capacitors_5_1/capacitor_5_4/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.98f
C624 cp2_buffer_5stage_0/cp2_buffer1_0/charge_pump_0/capacitors_5_1/capacitor_5_4/buffer_digital_1/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.58f
C625 cp2_buffer_5stage_0/cp2_buffer1_0/charge_pump_0/capacitors_5_1/capacitor_5_3/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.34f
C626 cp2_buffer_5stage_0/cp2_buffer1_0/charge_pump_0/capacitors_5_1/capacitor_5_3/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.98f
C627 cp2_buffer_5stage_0/cp2_buffer1_0/charge_pump_0/capacitors_5_1/capacitor_5_3/buffer_digital_1/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.58f
C628 cp2_buffer_5stage_0/cp2_buffer1_0/charge_pump_0/capacitors_5_1/capacitor_5_2/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.34f
C629 cp2_buffer_5stage_0/cp2_buffer1_0/charge_pump_0/capacitors_5_1/capacitor_5_2/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.98f
C630 cp2_buffer_5stage_0/cp2_buffer1_0/charge_pump_0/capacitors_5_1/capacitor_5_2/buffer_digital_1/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.58f
C631 cp2_buffer_5stage_0/cp2_buffer1_0/charge_pump_0/capacitors_5_1/capacitor_5_1/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.34f
C632 cp2_buffer_5stage_0/cp2_buffer1_0/charge_pump_0/capacitors_5_1/capacitor_5_1/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.98f
C633 cp2_buffer_5stage_0/cp2_buffer1_0/charge_pump_0/capacitors_5_1/capacitor_5_1/buffer_digital_1/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.58f
C634 cp2_buffer_5stage_0/cp2_buffer1_0/charge_pump_0/capacitors_5_1/capacitor_5_0/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.34f
C635 cp2_buffer_5stage_0/cp2_buffer1_0/charge_pump_0/capacitors_5_1/capacitor_5_0/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.98f
C636 cp2_buffer_5stage_0/cp2_buffer1_0/charge_pump_0/capacitors_5_1/capacitor_5_0/buffer_digital_1/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.58f
C637 cp2_buffer_5stage_0/cp2_buffer1_0/charge_pump_0/input2 cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 14.4f
C638 cp2_buffer_5stage_0/cp2_buffer1_0/charge_pump_0/capacitors_5_1/capacitor_5_7/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.34f
C639 cp2_buffer_5stage_0/cp2_buffer1_0/charge_pump_0/clkb cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 84f
C640 cp2_buffer_5stage_0/cp2_buffer1_0/charge_pump_0/capacitors_5_1/capacitor_5_7/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.98f
C641 cp2_buffer_5stage_0/cp2_buffer1_0/charge_pump_0/capacitors_5_1/capacitor_5_7/buffer_digital_1/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.58f
C642 cp2_buffer_5stage_0/cp2_buffer1_0/charge_pump_0/capacitors_5_1/capacitor_5_6/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.34f
C643 cp2_buffer_5stage_0/cp2_buffer1_0/charge_pump_0/capacitors_5_1/capacitor_5_6/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.98f
C644 cp2_buffer_5stage_0/cp2_buffer1_0/charge_pump_0/capacitors_5_1/capacitor_5_6/buffer_digital_1/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.58f
C645 cp2_buffer_5stage_0/cp2_buffer1_0/charge_pump_0/capacitors_5_1/capacitor_5_5/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.34f
C646 cp2_buffer_5stage_0/cp2_buffer1_0/charge_pump_0/capacitors_5_1/capacitor_5_5/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.98f
C647 cp2_buffer_5stage_0/cp2_buffer1_0/charge_pump_0/capacitors_5_1/capacitor_5_5/buffer_digital_1/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.58f
C648 cp2_buffer_5stage_0/cp2_buffer1_0/charge_pump_0/g1 cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.63f
C649 cp1_buffer_5stage_0/cp1_buffer1_reverse_1/charge_pump1_reverse_0/input1 cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 22.6f
C650 cp1_buffer_5stage_0/cp1_buffer1_reverse_1/charge_pump1_reverse_0/capacitors_1_12/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.34f
C651 cp1_buffer_5stage_0/cp1_buffer1_reverse_1/charge_pump1_reverse_0/capacitors_1_12/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.98f
C652 cp1_buffer_5stage_0/cp1_buffer1_reverse_1/charge_pump1_reverse_0/capacitors_1_12/capacitor_8_0/capacitor_7_0/buffer_digital_0/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.61f
C653 cp1_buffer_5stage_0/cp1_buffer1_reverse_1/charge_pump1_reverse_0/capacitors_1_13/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.34f
C654 cp1_buffer_5stage_0/cp1_buffer1_reverse_1/charge_pump1_reverse_0/capacitors_1_13/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.98f
C655 cp1_buffer_5stage_0/cp1_buffer1_reverse_1/charge_pump1_reverse_0/capacitors_1_13/capacitor_8_0/capacitor_7_0/buffer_digital_0/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.61f
C656 cp1_buffer_5stage_0/cp1_buffer1_reverse_1/charge_pump1_reverse_0/capacitors_1_11/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.34f
C657 cp1_buffer_5stage_0/cp1_buffer1_reverse_1/charge_pump1_reverse_0/capacitors_1_11/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.98f
C658 cp1_buffer_5stage_0/cp1_buffer1_reverse_1/charge_pump1_reverse_0/capacitors_1_11/capacitor_8_0/capacitor_7_0/buffer_digital_0/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.61f
C659 cp1_buffer_5stage_0/cp1_buffer1_reverse_1/charge_pump1_reverse_0/capacitors_1_10/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.34f
C660 cp1_buffer_5stage_0/cp1_buffer1_reverse_1/charge_pump1_reverse_0/capacitors_1_10/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.98f
C661 cp1_buffer_5stage_0/cp1_buffer1_reverse_1/charge_pump1_reverse_0/capacitors_1_10/capacitor_8_0/capacitor_7_0/buffer_digital_0/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.61f
C662 cp1_buffer_5stage_0/cp1_buffer1_reverse_1/charge_pump1_reverse_0/m1_4341_n519# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 3.33f
C663 cp1_buffer_5stage_0/cp1_buffer1_reverse_1/charge_pump1_reverse_0/input2 cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 22.2f
C664 cp1_buffer_5stage_0/cp1_buffer1_reverse_1/charge_pump1_reverse_0/m1_12659_300# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.68f
C665 cp1_buffer_5stage_0/cp1_buffer1_reverse_1/charge_pump1_reverse_0/capacitors_1_9/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.34f
C666 cp1_buffer_5stage_0/cp1_buffer1_reverse_1/charge_pump1_reverse_0/capacitors_1_9/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.98f
C667 cp1_buffer_5stage_0/cp1_buffer1_reverse_1/charge_pump1_reverse_0/capacitors_1_9/capacitor_8_0/capacitor_7_0/buffer_digital_0/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.61f
C668 cp1_buffer_5stage_0/cp1_buffer1_reverse_1/charge_pump1_reverse_0/capacitors_1_8/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.34f
C669 cp1_buffer_5stage_0/cp1_buffer1_reverse_1/charge_pump1_reverse_0/capacitors_1_8/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.98f
C670 cp1_buffer_5stage_0/cp1_buffer1_reverse_1/charge_pump1_reverse_0/capacitors_1_8/capacitor_8_0/capacitor_7_0/buffer_digital_0/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.61f
C671 cp1_buffer_5stage_0/cp1_buffer1_reverse_1/charge_pump1_reverse_0/capacitors_1_7/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.34f
C672 cp1_buffer_5stage_0/cp1_buffer1_reverse_1/charge_pump1_reverse_0/capacitors_1_7/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.98f
C673 cp1_buffer_5stage_0/cp1_buffer1_reverse_1/charge_pump1_reverse_0/capacitors_1_7/capacitor_8_0/capacitor_7_0/buffer_digital_0/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.61f
C674 cp1_buffer_5stage_0/cp1_buffer1_reverse_1/charge_pump1_reverse_0/capacitors_1_6/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.34f
C675 cp1_buffer_5stage_0/cp1_buffer1_reverse_1/charge_pump1_reverse_0/capacitors_1_6/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.98f
C676 cp1_buffer_5stage_0/cp1_buffer1_reverse_1/charge_pump1_reverse_0/capacitors_1_6/capacitor_8_0/capacitor_7_0/buffer_digital_0/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.61f
C677 cp1_buffer_5stage_0/cp1_buffer1_reverse_1/charge_pump1_reverse_0/capacitors_1_5/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.34f
C678 cp1_buffer_5stage_0/cp1_buffer1_reverse_1/charge_pump1_reverse_0/capacitors_1_5/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.98f
C679 cp1_buffer_5stage_0/cp1_buffer1_reverse_1/charge_pump1_reverse_0/capacitors_1_5/capacitor_8_0/capacitor_7_0/buffer_digital_0/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.61f
C680 cp1_buffer_5stage_0/cp1_buffer1_reverse_1/charge_pump1_reverse_0/capacitors_1_4/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.34f
C681 cp1_buffer_5stage_0/cp1_buffer1_reverse_1/charge_pump1_reverse_0/capacitors_1_4/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.98f
C682 cp1_buffer_5stage_0/cp1_buffer1_reverse_1/charge_pump1_reverse_0/capacitors_1_4/capacitor_8_0/capacitor_7_0/buffer_digital_0/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.61f
C683 cp1_buffer_5stage_0/cp1_buffer1_reverse_1/charge_pump1_reverse_0/capacitors_1_3/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.34f
C684 cp1_buffer_5stage_0/cp1_buffer1_reverse_1/charge_pump1_reverse_0/capacitors_1_3/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.98f
C685 cp1_buffer_5stage_0/cp1_buffer1_reverse_1/charge_pump1_reverse_0/capacitors_1_3/capacitor_8_0/capacitor_7_0/buffer_digital_0/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.61f
C686 cp1_buffer_5stage_0/cp1_buffer1_reverse_1/charge_pump1_reverse_0/capacitors_1_2/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.34f
C687 cp1_buffer_5stage_0/cp1_buffer1_reverse_1/charge_pump1_reverse_0/capacitors_1_2/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.98f
C688 cp1_buffer_5stage_0/cp1_buffer1_reverse_1/charge_pump1_reverse_0/capacitors_1_2/capacitor_8_0/capacitor_7_0/buffer_digital_0/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.61f
C689 cp1_buffer_5stage_0/cp1_buffer1_reverse_1/charge_pump1_reverse_0/capacitors_1_1/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.34f
C690 cp1_buffer_5stage_0/cp1_buffer1_reverse_1/charge_pump1_reverse_0/capacitors_1_1/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.98f
C691 cp1_buffer_5stage_0/cp1_buffer1_reverse_1/charge_pump1_reverse_0/capacitors_1_1/capacitor_8_0/capacitor_7_0/buffer_digital_0/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.61f
C692 cp1_buffer_5stage_0/cp1_buffer1_reverse_1/charge_pump1_reverse_0/capacitors_1_0/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.34f
C693 cp1_buffer_5stage_0/cp1_buffer1_reverse_1/charge_pump1_reverse_0/capacitors_1_0/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.98f
C694 cp1_buffer_5stage_0/cp1_buffer1_reverse_1/charge_pump1_reverse_0/capacitors_1_0/capacitor_8_0/capacitor_7_0/buffer_digital_0/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.61f
C695 cp1_buffer_5stage_0/cp1_buffer1_reverse_1/charge_pump1_reverse_0/capacitor_8_1/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.34f
C696 cp1_buffer_5stage_0/cp1_buffer1_reverse_1/charge_pump1_reverse_0/clock_1/clk cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 94.6f
C697 cp1_buffer_5stage_0/cp1_buffer1_reverse_1/charge_pump1_reverse_0/capacitor_8_1/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.98f
C698 cp1_buffer_5stage_0/cp1_buffer1_reverse_1/charge_pump1_reverse_0/capacitor_8_1/capacitor_7_0/buffer_digital_0/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.61f
C699 cp1_buffer_5stage_0/cp1_buffer1_reverse_1/charge_pump1_reverse_0/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.34f
C700 cp1_buffer_5stage_0/cp1_buffer1_reverse_1/charge_pump1_reverse_0/clock_1/clkb cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 0.101p
C701 cp1_buffer_5stage_0/cp1_buffer1_reverse_1/charge_pump1_reverse_0/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.98f
C702 cp1_buffer_5stage_0/cp1_buffer1_reverse_1/charge_pump1_reverse_0/capacitor_8_0/capacitor_7_0/buffer_digital_0/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.61f
C703 cp1_buffer_5stage_0/cp1_buffer1_reverse_1/charge_pump1_reverse_0/clock_1/a_2432_n962# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 8.68f **FLOATING
C704 cp1_buffer_5stage_0/cp1_buffer1_reverse_1/charge_pump1_reverse_0/clock_1/a_2020_n482# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.57f **FLOATING
C705 cp1_buffer_5stage_0/cp1_buffer1_reverse_1/charge_pump1_reverse_0/clock_1/a_344_102# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.81f
C706 cp1_buffer_5stage_0/cp1_buffer1_reverse_1/charge_pump1_reverse_0/clock_1/a_2402_572# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.17f
C707 cp1_buffer_5stage_0/cp1_buffer1_reverse_1/charge_pump1_reverse_0/clock_1/a_344_n986# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.38f
C708 cp1_buffer_5stage_0/cp1_buffer1_2/clk_in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 5.35f
C709 cp1_buffer_5stage_0/cp1_buffer1_reverse_1/charge_pump1_reverse_0/clock_1/a_3246_118# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 6.83f
C710 cp1_buffer_5stage_0/cp1_buffer1_reverse_0/charge_pump1_reverse_0/input1 cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 22.6f
C711 cp1_buffer_5stage_0/cp1_buffer1_reverse_0/charge_pump1_reverse_0/capacitors_1_12/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.34f
C712 cp1_buffer_5stage_0/cp1_buffer1_reverse_0/charge_pump1_reverse_0/capacitors_1_12/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.98f
C713 cp1_buffer_5stage_0/cp1_buffer1_reverse_0/charge_pump1_reverse_0/capacitors_1_12/capacitor_8_0/capacitor_7_0/buffer_digital_0/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.61f
C714 cp1_buffer_5stage_0/cp1_buffer1_reverse_0/charge_pump1_reverse_0/capacitors_1_13/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.34f
C715 cp1_buffer_5stage_0/cp1_buffer1_reverse_0/charge_pump1_reverse_0/capacitors_1_13/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.98f
C716 cp1_buffer_5stage_0/cp1_buffer1_reverse_0/charge_pump1_reverse_0/capacitors_1_13/capacitor_8_0/capacitor_7_0/buffer_digital_0/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.61f
C717 cp1_buffer_5stage_0/cp1_buffer1_reverse_0/charge_pump1_reverse_0/capacitors_1_11/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.34f
C718 cp1_buffer_5stage_0/cp1_buffer1_reverse_0/charge_pump1_reverse_0/capacitors_1_11/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.98f
C719 cp1_buffer_5stage_0/cp1_buffer1_reverse_0/charge_pump1_reverse_0/capacitors_1_11/capacitor_8_0/capacitor_7_0/buffer_digital_0/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.61f
C720 cp1_buffer_5stage_0/cp1_buffer1_reverse_0/charge_pump1_reverse_0/capacitors_1_10/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.34f
C721 cp1_buffer_5stage_0/cp1_buffer1_reverse_0/charge_pump1_reverse_0/capacitors_1_10/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.98f
C722 cp1_buffer_5stage_0/cp1_buffer1_reverse_0/charge_pump1_reverse_0/capacitors_1_10/capacitor_8_0/capacitor_7_0/buffer_digital_0/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.61f
C723 cp1_buffer_5stage_0/cp1_buffer1_reverse_0/charge_pump1_reverse_0/m1_4341_n519# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 3.33f
C724 cp1_buffer_5stage_0/cp1_buffer1_reverse_0/charge_pump1_reverse_0/input2 cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 22.2f
C725 cp1_buffer_5stage_0/cp1_buffer1_reverse_0/charge_pump1_reverse_0/m1_12659_300# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.68f
C726 cp1_buffer_5stage_0/cp1_buffer1_reverse_0/charge_pump1_reverse_0/capacitors_1_9/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.34f
C727 cp1_buffer_5stage_0/cp1_buffer1_reverse_0/charge_pump1_reverse_0/capacitors_1_9/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.98f
C728 cp1_buffer_5stage_0/cp1_buffer1_reverse_0/charge_pump1_reverse_0/capacitors_1_9/capacitor_8_0/capacitor_7_0/buffer_digital_0/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.61f
C729 cp1_buffer_5stage_0/cp1_buffer1_reverse_0/charge_pump1_reverse_0/capacitors_1_8/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.34f
C730 cp1_buffer_5stage_0/cp1_buffer1_reverse_0/charge_pump1_reverse_0/capacitors_1_8/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.98f
C731 cp1_buffer_5stage_0/cp1_buffer1_reverse_0/charge_pump1_reverse_0/capacitors_1_8/capacitor_8_0/capacitor_7_0/buffer_digital_0/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.61f
C732 cp1_buffer_5stage_0/cp1_buffer1_reverse_0/charge_pump1_reverse_0/capacitors_1_7/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.34f
C733 cp1_buffer_5stage_0/cp1_buffer1_reverse_0/charge_pump1_reverse_0/capacitors_1_7/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.98f
C734 cp1_buffer_5stage_0/cp1_buffer1_reverse_0/charge_pump1_reverse_0/capacitors_1_7/capacitor_8_0/capacitor_7_0/buffer_digital_0/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.61f
C735 cp1_buffer_5stage_0/cp1_buffer1_reverse_0/charge_pump1_reverse_0/capacitors_1_6/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.34f
C736 cp1_buffer_5stage_0/cp1_buffer1_reverse_0/charge_pump1_reverse_0/capacitors_1_6/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.98f
C737 cp1_buffer_5stage_0/cp1_buffer1_reverse_0/charge_pump1_reverse_0/capacitors_1_6/capacitor_8_0/capacitor_7_0/buffer_digital_0/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.61f
C738 cp1_buffer_5stage_0/cp1_buffer1_reverse_0/charge_pump1_reverse_0/capacitors_1_5/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.34f
C739 cp1_buffer_5stage_0/cp1_buffer1_reverse_0/charge_pump1_reverse_0/capacitors_1_5/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.98f
C740 cp1_buffer_5stage_0/cp1_buffer1_reverse_0/charge_pump1_reverse_0/capacitors_1_5/capacitor_8_0/capacitor_7_0/buffer_digital_0/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.61f
C741 cp1_buffer_5stage_0/cp1_buffer1_reverse_0/charge_pump1_reverse_0/capacitors_1_4/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.34f
C742 cp1_buffer_5stage_0/cp1_buffer1_reverse_0/charge_pump1_reverse_0/capacitors_1_4/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.98f
C743 cp1_buffer_5stage_0/cp1_buffer1_reverse_0/charge_pump1_reverse_0/capacitors_1_4/capacitor_8_0/capacitor_7_0/buffer_digital_0/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.61f
C744 cp1_buffer_5stage_0/cp1_buffer1_reverse_0/charge_pump1_reverse_0/capacitors_1_3/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.34f
C745 cp1_buffer_5stage_0/cp1_buffer1_reverse_0/charge_pump1_reverse_0/capacitors_1_3/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.98f
C746 cp1_buffer_5stage_0/cp1_buffer1_reverse_0/charge_pump1_reverse_0/capacitors_1_3/capacitor_8_0/capacitor_7_0/buffer_digital_0/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.61f
C747 cp1_buffer_5stage_0/cp1_buffer1_reverse_0/charge_pump1_reverse_0/capacitors_1_2/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.34f
C748 cp1_buffer_5stage_0/cp1_buffer1_reverse_0/charge_pump1_reverse_0/capacitors_1_2/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.98f
C749 cp1_buffer_5stage_0/cp1_buffer1_reverse_0/charge_pump1_reverse_0/capacitors_1_2/capacitor_8_0/capacitor_7_0/buffer_digital_0/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.61f
C750 cp1_buffer_5stage_0/cp1_buffer1_reverse_0/charge_pump1_reverse_0/capacitors_1_1/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.34f
C751 cp1_buffer_5stage_0/cp1_buffer1_reverse_0/charge_pump1_reverse_0/capacitors_1_1/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.98f
C752 cp1_buffer_5stage_0/cp1_buffer1_reverse_0/charge_pump1_reverse_0/capacitors_1_1/capacitor_8_0/capacitor_7_0/buffer_digital_0/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.61f
C753 cp1_buffer_5stage_0/cp1_buffer1_reverse_0/charge_pump1_reverse_0/capacitors_1_0/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.34f
C754 cp1_buffer_5stage_0/cp1_buffer1_reverse_0/charge_pump1_reverse_0/capacitors_1_0/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.98f
C755 cp1_buffer_5stage_0/cp1_buffer1_reverse_0/charge_pump1_reverse_0/capacitors_1_0/capacitor_8_0/capacitor_7_0/buffer_digital_0/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.61f
C756 cp1_buffer_5stage_0/cp1_buffer1_reverse_0/charge_pump1_reverse_0/capacitor_8_1/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.34f
C757 cp1_buffer_5stage_0/cp1_buffer1_reverse_0/charge_pump1_reverse_0/clock_1/clk cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 94.6f
C758 cp1_buffer_5stage_0/cp1_buffer1_reverse_0/charge_pump1_reverse_0/capacitor_8_1/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.98f
C759 cp1_buffer_5stage_0/cp1_buffer1_reverse_0/charge_pump1_reverse_0/capacitor_8_1/capacitor_7_0/buffer_digital_0/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.61f
C760 cp1_buffer_5stage_0/cp1_buffer1_reverse_0/charge_pump1_reverse_0/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.34f
C761 cp1_buffer_5stage_0/cp1_buffer1_reverse_0/charge_pump1_reverse_0/clock_1/clkb cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 0.101p
C762 cp1_buffer_5stage_0/cp1_buffer1_reverse_0/charge_pump1_reverse_0/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.98f
C763 cp1_buffer_5stage_0/cp1_buffer1_reverse_0/charge_pump1_reverse_0/capacitor_8_0/capacitor_7_0/buffer_digital_0/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.61f
C764 cp1_buffer_5stage_0/cp1_buffer1_reverse_0/charge_pump1_reverse_0/clock_1/a_2432_n962# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 8.68f **FLOATING
C765 cp1_buffer_5stage_0/cp1_buffer1_reverse_0/charge_pump1_reverse_0/clock_1/a_2020_n482# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.57f **FLOATING
C766 cp1_buffer_5stage_0/cp1_buffer1_reverse_0/charge_pump1_reverse_0/clock_1/a_344_102# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.81f
C767 cp1_buffer_5stage_0/cp1_buffer1_reverse_0/charge_pump1_reverse_0/clock_1/a_2402_572# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.17f
C768 cp1_buffer_5stage_0/cp1_buffer1_reverse_0/charge_pump1_reverse_0/clock_1/a_344_n986# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.38f
C769 cp1_buffer_5stage_0/cp1_buffer1_1/clk_in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 4.43f
C770 cp1_buffer_5stage_0/cp1_buffer1_reverse_0/charge_pump1_reverse_0/clock_1/a_3246_118# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 6.83f
C771 cp1_buffer_5stage_0/cp1_buffer1_2/clk_out cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 3.51f
C772 cp1_buffer_5stage_0/cp1_buffer1_2/charge_pump1_0/input1 cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 22.5f
C773 cp1_buffer_5stage_0/cp1_buffer1_2/charge_pump1_0/input2 cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 22.2f
C774 cp1_buffer_5stage_0/cp1_buffer1_2/charge_pump1_0/capacitors_1_12/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.34f
C775 cp1_buffer_5stage_0/cp1_buffer1_2/charge_pump1_0/capacitors_1_12/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.98f
C776 cp1_buffer_5stage_0/cp1_buffer1_2/charge_pump1_0/capacitors_1_12/capacitor_8_0/capacitor_7_0/buffer_digital_0/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.61f
C777 cp1_buffer_5stage_0/cp1_buffer1_2/charge_pump1_0/capacitors_1_13/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.34f
C778 cp1_buffer_5stage_0/cp1_buffer1_2/charge_pump1_0/capacitors_1_13/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.98f
C779 cp1_buffer_5stage_0/cp1_buffer1_2/charge_pump1_0/capacitors_1_13/capacitor_8_0/capacitor_7_0/buffer_digital_0/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.61f
C780 cp1_buffer_5stage_0/cp1_buffer1_2/charge_pump1_0/capacitors_1_11/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.34f
C781 cp1_buffer_5stage_0/cp1_buffer1_2/charge_pump1_0/capacitors_1_11/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.98f
C782 cp1_buffer_5stage_0/cp1_buffer1_2/charge_pump1_0/capacitors_1_11/capacitor_8_0/capacitor_7_0/buffer_digital_0/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.61f
C783 cp1_buffer_5stage_0/cp1_buffer1_2/charge_pump1_0/capacitors_1_10/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.34f
C784 cp1_buffer_5stage_0/cp1_buffer1_2/charge_pump1_0/capacitors_1_10/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.98f
C785 cp1_buffer_5stage_0/cp1_buffer1_2/charge_pump1_0/capacitors_1_10/capacitor_8_0/capacitor_7_0/buffer_digital_0/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.61f
C786 cp1_buffer_5stage_0/cp1_buffer1_2/charge_pump1_0/m1_4341_n519# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 3.77f
C787 cp1_buffer_5stage_0/cp1_buffer1_2/charge_pump1_0/m1_12659_300# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.54f
C788 cp1_buffer_5stage_0/cp1_buffer1_2/charge_pump1_0/capacitors_1_9/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.34f
C789 cp1_buffer_5stage_0/cp1_buffer1_2/charge_pump1_0/capacitors_1_9/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.98f
C790 cp1_buffer_5stage_0/cp1_buffer1_2/charge_pump1_0/capacitors_1_9/capacitor_8_0/capacitor_7_0/buffer_digital_0/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.61f
C791 cp1_buffer_5stage_0/cp1_buffer1_2/charge_pump1_0/capacitors_1_8/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.34f
C792 cp1_buffer_5stage_0/cp1_buffer1_2/charge_pump1_0/capacitors_1_8/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.98f
C793 cp1_buffer_5stage_0/cp1_buffer1_2/charge_pump1_0/capacitors_1_8/capacitor_8_0/capacitor_7_0/buffer_digital_0/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.61f
C794 cp1_buffer_5stage_0/cp1_buffer1_2/charge_pump1_0/capacitors_1_7/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.34f
C795 cp1_buffer_5stage_0/cp1_buffer1_2/charge_pump1_0/capacitors_1_7/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.98f
C796 cp1_buffer_5stage_0/cp1_buffer1_2/charge_pump1_0/capacitors_1_7/capacitor_8_0/capacitor_7_0/buffer_digital_0/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.61f
C797 cp1_buffer_5stage_0/cp1_buffer1_2/charge_pump1_0/capacitors_1_6/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.34f
C798 cp1_buffer_5stage_0/cp1_buffer1_2/charge_pump1_0/capacitors_1_6/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.98f
C799 cp1_buffer_5stage_0/cp1_buffer1_2/charge_pump1_0/capacitors_1_6/capacitor_8_0/capacitor_7_0/buffer_digital_0/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.61f
C800 cp1_buffer_5stage_0/cp1_buffer1_2/charge_pump1_0/capacitors_1_5/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.34f
C801 cp1_buffer_5stage_0/cp1_buffer1_2/charge_pump1_0/capacitors_1_5/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.98f
C802 cp1_buffer_5stage_0/cp1_buffer1_2/charge_pump1_0/capacitors_1_5/capacitor_8_0/capacitor_7_0/buffer_digital_0/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.61f
C803 cp1_buffer_5stage_0/cp1_buffer1_2/charge_pump1_0/capacitors_1_4/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.34f
C804 cp1_buffer_5stage_0/cp1_buffer1_2/charge_pump1_0/capacitors_1_4/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.98f
C805 cp1_buffer_5stage_0/cp1_buffer1_2/charge_pump1_0/capacitors_1_4/capacitor_8_0/capacitor_7_0/buffer_digital_0/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.61f
C806 cp1_buffer_5stage_0/cp1_buffer1_2/charge_pump1_0/capacitors_1_3/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.34f
C807 cp1_buffer_5stage_0/cp1_buffer1_2/charge_pump1_0/capacitors_1_3/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.98f
C808 cp1_buffer_5stage_0/cp1_buffer1_2/charge_pump1_0/capacitors_1_3/capacitor_8_0/capacitor_7_0/buffer_digital_0/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.61f
C809 cp1_buffer_5stage_0/cp1_buffer1_2/charge_pump1_0/capacitors_1_2/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.34f
C810 cp1_buffer_5stage_0/cp1_buffer1_2/charge_pump1_0/capacitors_1_2/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.98f
C811 cp1_buffer_5stage_0/cp1_buffer1_2/charge_pump1_0/capacitors_1_2/capacitor_8_0/capacitor_7_0/buffer_digital_0/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.61f
C812 cp1_buffer_5stage_0/cp1_buffer1_2/charge_pump1_0/capacitors_1_1/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.34f
C813 cp1_buffer_5stage_0/cp1_buffer1_2/charge_pump1_0/capacitors_1_1/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.98f
C814 cp1_buffer_5stage_0/cp1_buffer1_2/charge_pump1_0/capacitors_1_1/capacitor_8_0/capacitor_7_0/buffer_digital_0/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.61f
C815 cp1_buffer_5stage_0/cp1_buffer1_2/charge_pump1_0/capacitors_1_0/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.34f
C816 cp1_buffer_5stage_0/cp1_buffer1_2/charge_pump1_0/capacitors_1_0/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.98f
C817 cp1_buffer_5stage_0/cp1_buffer1_2/charge_pump1_0/capacitors_1_0/capacitor_8_0/capacitor_7_0/buffer_digital_0/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.61f
C818 cp1_buffer_5stage_0/cp1_buffer1_2/charge_pump1_0/capacitor_8_1/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.34f
C819 cp1_buffer_5stage_0/cp1_buffer1_2/charge_pump1_0/clkb cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 89.9f
C820 cp1_buffer_5stage_0/cp1_buffer1_2/charge_pump1_0/capacitor_8_1/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.98f
C821 cp1_buffer_5stage_0/cp1_buffer1_2/charge_pump1_0/capacitor_8_1/capacitor_7_0/buffer_digital_0/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.61f
C822 cp1_buffer_5stage_0/cp1_buffer1_2/charge_pump1_0/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.34f
C823 cp1_buffer_5stage_0/cp1_buffer1_2/charge_pump1_0/clk cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 89f
C824 cp1_buffer_5stage_0/cp1_buffer1_2/charge_pump1_0/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.98f
C825 cp1_buffer_5stage_0/cp1_buffer1_2/charge_pump1_0/capacitor_8_0/capacitor_7_0/buffer_digital_0/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.61f
C826 cp1_buffer_5stage_0/cp1_buffer1_2/charge_pump1_0/clock_0/a_2432_n962# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 8.68f **FLOATING
C827 cp1_buffer_5stage_0/cp1_buffer1_2/charge_pump1_0/clock_0/a_2020_n482# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.57f **FLOATING
C828 cp1_buffer_5stage_0/cp1_buffer1_2/charge_pump1_0/clock_0/a_344_102# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.81f
C829 cp1_buffer_5stage_0/cp1_buffer1_2/charge_pump1_0/clock_0/a_2402_572# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.17f
C830 cp1_buffer_5stage_0/cp1_buffer1_2/charge_pump1_0/clock_0/a_344_n986# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.38f
C831 cp1_buffer_5stage_0/cp1_buffer1_2/charge_pump1_0/clock_0/a_3246_118# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 6.83f
C832 cp1_buffer_5stage_0/cp1_buffer1_2/charge_pump1_0/g2 cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.34f
C833 cp2_buffer_5stage_0/cp2_buffer1_0/charge_pump_0/vs cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 40.1f
C834 cp1_buffer_5stage_0/cp1_buffer1_1/clk_out cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 7.47f
C835 cp1_buffer_5stage_0/cp1_buffer1_1/charge_pump1_0/input1 cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 22.5f
C836 cp1_buffer_5stage_0/cp1_buffer1_1/charge_pump1_0/input2 cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 22.2f
C837 cp1_buffer_5stage_0/cp1_buffer1_1/charge_pump1_0/capacitors_1_12/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.34f
C838 cp1_buffer_5stage_0/cp1_buffer1_1/charge_pump1_0/capacitors_1_12/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.98f
C839 cp1_buffer_5stage_0/cp1_buffer1_1/charge_pump1_0/capacitors_1_12/capacitor_8_0/capacitor_7_0/buffer_digital_0/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.61f
C840 cp1_buffer_5stage_0/cp1_buffer1_1/charge_pump1_0/capacitors_1_13/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.34f
C841 cp1_buffer_5stage_0/cp1_buffer1_1/charge_pump1_0/capacitors_1_13/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.98f
C842 cp1_buffer_5stage_0/cp1_buffer1_1/charge_pump1_0/capacitors_1_13/capacitor_8_0/capacitor_7_0/buffer_digital_0/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.61f
C843 cp1_buffer_5stage_0/cp1_buffer1_1/charge_pump1_0/capacitors_1_11/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.34f
C844 cp1_buffer_5stage_0/cp1_buffer1_1/charge_pump1_0/capacitors_1_11/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.98f
C845 cp1_buffer_5stage_0/cp1_buffer1_1/charge_pump1_0/capacitors_1_11/capacitor_8_0/capacitor_7_0/buffer_digital_0/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.61f
C846 cp1_buffer_5stage_0/cp1_buffer1_1/charge_pump1_0/capacitors_1_10/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.34f
C847 cp1_buffer_5stage_0/cp1_buffer1_1/charge_pump1_0/capacitors_1_10/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.98f
C848 cp1_buffer_5stage_0/cp1_buffer1_1/charge_pump1_0/capacitors_1_10/capacitor_8_0/capacitor_7_0/buffer_digital_0/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.61f
C849 cp1_buffer_5stage_0/cp1_buffer1_1/charge_pump1_0/m1_4341_n519# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 3.77f
C850 cp1_buffer_5stage_0/cp1_buffer1_1/charge_pump1_0/m1_12659_300# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.54f
C851 cp1_buffer_5stage_0/cp1_buffer1_reverse_1/charge_pump1_reverse_0/nmos_dnw3_0/vs cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 14.5f
C852 cp1_buffer_5stage_0/cp1_buffer1_1/charge_pump1_0/capacitors_1_9/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.34f
C853 cp1_buffer_5stage_0/cp1_buffer1_1/charge_pump1_0/capacitors_1_9/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.98f
C854 cp1_buffer_5stage_0/cp1_buffer1_1/charge_pump1_0/capacitors_1_9/capacitor_8_0/capacitor_7_0/buffer_digital_0/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.61f
C855 cp1_buffer_5stage_0/cp1_buffer1_1/charge_pump1_0/capacitors_1_8/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.34f
C856 cp1_buffer_5stage_0/cp1_buffer1_1/charge_pump1_0/capacitors_1_8/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.98f
C857 cp1_buffer_5stage_0/cp1_buffer1_1/charge_pump1_0/capacitors_1_8/capacitor_8_0/capacitor_7_0/buffer_digital_0/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.61f
C858 cp1_buffer_5stage_0/cp1_buffer1_1/charge_pump1_0/capacitors_1_7/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.34f
C859 cp1_buffer_5stage_0/cp1_buffer1_1/charge_pump1_0/capacitors_1_7/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.98f
C860 cp1_buffer_5stage_0/cp1_buffer1_1/charge_pump1_0/capacitors_1_7/capacitor_8_0/capacitor_7_0/buffer_digital_0/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.61f
C861 cp1_buffer_5stage_0/cp1_buffer1_1/charge_pump1_0/capacitors_1_6/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.34f
C862 cp1_buffer_5stage_0/cp1_buffer1_1/charge_pump1_0/capacitors_1_6/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.98f
C863 cp1_buffer_5stage_0/cp1_buffer1_1/charge_pump1_0/capacitors_1_6/capacitor_8_0/capacitor_7_0/buffer_digital_0/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.61f
C864 cp1_buffer_5stage_0/cp1_buffer1_1/charge_pump1_0/capacitors_1_5/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.34f
C865 cp1_buffer_5stage_0/cp1_buffer1_1/charge_pump1_0/capacitors_1_5/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.98f
C866 cp1_buffer_5stage_0/cp1_buffer1_1/charge_pump1_0/capacitors_1_5/capacitor_8_0/capacitor_7_0/buffer_digital_0/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.61f
C867 cp1_buffer_5stage_0/cp1_buffer1_1/charge_pump1_0/capacitors_1_4/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.34f
C868 cp1_buffer_5stage_0/cp1_buffer1_1/charge_pump1_0/capacitors_1_4/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.98f
C869 cp1_buffer_5stage_0/cp1_buffer1_1/charge_pump1_0/capacitors_1_4/capacitor_8_0/capacitor_7_0/buffer_digital_0/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.61f
C870 cp1_buffer_5stage_0/cp1_buffer1_1/charge_pump1_0/capacitors_1_3/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.34f
C871 cp1_buffer_5stage_0/cp1_buffer1_1/charge_pump1_0/capacitors_1_3/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.98f
C872 cp1_buffer_5stage_0/cp1_buffer1_1/charge_pump1_0/capacitors_1_3/capacitor_8_0/capacitor_7_0/buffer_digital_0/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.61f
C873 cp1_buffer_5stage_0/cp1_buffer1_1/charge_pump1_0/capacitors_1_2/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.34f
C874 cp1_buffer_5stage_0/cp1_buffer1_1/charge_pump1_0/capacitors_1_2/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.98f
C875 cp1_buffer_5stage_0/cp1_buffer1_1/charge_pump1_0/capacitors_1_2/capacitor_8_0/capacitor_7_0/buffer_digital_0/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.61f
C876 cp1_buffer_5stage_0/cp1_buffer1_1/charge_pump1_0/capacitors_1_1/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.34f
C877 cp1_buffer_5stage_0/cp1_buffer1_1/charge_pump1_0/capacitors_1_1/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.98f
C878 cp1_buffer_5stage_0/cp1_buffer1_1/charge_pump1_0/capacitors_1_1/capacitor_8_0/capacitor_7_0/buffer_digital_0/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.61f
C879 cp1_buffer_5stage_0/cp1_buffer1_1/charge_pump1_0/capacitors_1_0/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.34f
C880 cp1_buffer_5stage_0/cp1_buffer1_1/charge_pump1_0/capacitors_1_0/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.98f
C881 cp1_buffer_5stage_0/cp1_buffer1_1/charge_pump1_0/capacitors_1_0/capacitor_8_0/capacitor_7_0/buffer_digital_0/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.61f
C882 cp1_buffer_5stage_0/cp1_buffer1_1/charge_pump1_0/capacitor_8_1/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.34f
C883 cp1_buffer_5stage_0/cp1_buffer1_1/charge_pump1_0/clkb cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 89.9f
C884 cp1_buffer_5stage_0/cp1_buffer1_1/charge_pump1_0/capacitor_8_1/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.98f
C885 cp1_buffer_5stage_0/cp1_buffer1_1/charge_pump1_0/capacitor_8_1/capacitor_7_0/buffer_digital_0/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.61f
C886 cp1_buffer_5stage_0/cp1_buffer1_1/charge_pump1_0/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.34f
C887 cp1_buffer_5stage_0/cp1_buffer1_1/charge_pump1_0/clk cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 89f
C888 cp1_buffer_5stage_0/cp1_buffer1_1/charge_pump1_0/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.98f
C889 cp1_buffer_5stage_0/cp1_buffer1_1/charge_pump1_0/capacitor_8_0/capacitor_7_0/buffer_digital_0/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.61f
C890 cp1_buffer_5stage_0/cp1_buffer1_1/charge_pump1_0/clock_0/a_2432_n962# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 8.68f **FLOATING
C891 cp1_buffer_5stage_0/cp1_buffer1_1/charge_pump1_0/clock_0/a_2020_n482# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.57f **FLOATING
C892 cp1_buffer_5stage_0/cp1_buffer1_1/charge_pump1_0/clock_0/a_344_102# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.81f
C893 cp1_buffer_5stage_0/cp1_buffer1_1/charge_pump1_0/clock_0/a_2402_572# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.17f
C894 cp1_buffer_5stage_0/cp1_buffer1_1/charge_pump1_0/clock_0/a_344_n986# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.38f
C895 cp1_buffer_5stage_0/cp1_buffer1_1/charge_pump1_0/clock_0/a_3246_118# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 6.83f
C896 cp1_buffer_5stage_0/cp1_buffer1_1/charge_pump1_0/g2 cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.34f
C897 cp1_buffer_5stage_0/cp1_buffer1_1/charge_pump1_0/vin cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 13.2f
C898 cp1_buffer_5stage_0/cp1_buffer1_0/clk_in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 60.1f
C899 cp1_buffer_5stage_0/cp1_buffer1_0/clk_out cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 7.49f
C900 cp1_buffer_5stage_0/cp1_buffer1_0/charge_pump1_0/input1 cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 22.5f
C901 cp1_buffer_5stage_0/cp1_buffer1_0/charge_pump1_0/input2 cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 22.2f
C902 cp1_buffer_5stage_0/cp1_buffer1_0/charge_pump1_0/capacitors_1_12/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.34f
C903 cp1_buffer_5stage_0/cp1_buffer1_0/charge_pump1_0/capacitors_1_12/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.98f
C904 cp1_buffer_5stage_0/cp1_buffer1_0/charge_pump1_0/capacitors_1_12/capacitor_8_0/capacitor_7_0/buffer_digital_0/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.61f
C905 cp1_buffer_5stage_0/cp1_buffer1_0/charge_pump1_0/capacitors_1_13/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.34f
C906 cp1_buffer_5stage_0/cp1_buffer1_0/charge_pump1_0/capacitors_1_13/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.98f
C907 cp1_buffer_5stage_0/cp1_buffer1_0/charge_pump1_0/capacitors_1_13/capacitor_8_0/capacitor_7_0/buffer_digital_0/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.61f
C908 cp1_buffer_5stage_0/cp1_buffer1_0/charge_pump1_0/capacitors_1_11/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.34f
C909 cp1_buffer_5stage_0/cp1_buffer1_0/charge_pump1_0/capacitors_1_11/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.98f
C910 cp1_buffer_5stage_0/cp1_buffer1_0/charge_pump1_0/capacitors_1_11/capacitor_8_0/capacitor_7_0/buffer_digital_0/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.61f
C911 cp1_buffer_5stage_0/cp1_buffer1_0/charge_pump1_0/capacitors_1_10/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.34f
C912 cp1_buffer_5stage_0/cp1_buffer1_0/charge_pump1_0/capacitors_1_10/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.98f
C913 cp1_buffer_5stage_0/cp1_buffer1_0/charge_pump1_0/capacitors_1_10/capacitor_8_0/capacitor_7_0/buffer_digital_0/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.61f
C914 cp1_buffer_5stage_0/cp1_buffer1_0/charge_pump1_0/m1_4341_n519# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 3.77f
C915 cp1_buffer_5stage_0/cp1_buffer1_0/charge_pump1_0/m1_12659_300# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.54f
C916 cp1_buffer_5stage_0/cp1_buffer1_reverse_0/charge_pump1_reverse_0/nmos_dnw3_0/vs cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 14.6f
C917 cp1_buffer_5stage_0/cp1_buffer1_0/charge_pump1_0/capacitors_1_9/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.34f
C918 cp1_buffer_5stage_0/cp1_buffer1_0/charge_pump1_0/capacitors_1_9/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.98f
C919 cp1_buffer_5stage_0/cp1_buffer1_0/charge_pump1_0/capacitors_1_9/capacitor_8_0/capacitor_7_0/buffer_digital_0/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.61f
C920 cp1_buffer_5stage_0/cp1_buffer1_0/charge_pump1_0/capacitors_1_8/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.34f
C921 cp1_buffer_5stage_0/cp1_buffer1_0/charge_pump1_0/capacitors_1_8/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.98f
C922 cp1_buffer_5stage_0/cp1_buffer1_0/charge_pump1_0/capacitors_1_8/capacitor_8_0/capacitor_7_0/buffer_digital_0/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.61f
C923 cp1_buffer_5stage_0/cp1_buffer1_0/charge_pump1_0/capacitors_1_7/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.34f
C924 cp1_buffer_5stage_0/cp1_buffer1_0/charge_pump1_0/capacitors_1_7/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.98f
C925 cp1_buffer_5stage_0/cp1_buffer1_0/charge_pump1_0/capacitors_1_7/capacitor_8_0/capacitor_7_0/buffer_digital_0/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.61f
C926 cp1_buffer_5stage_0/cp1_buffer1_0/charge_pump1_0/capacitors_1_6/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.34f
C927 cp1_buffer_5stage_0/cp1_buffer1_0/charge_pump1_0/capacitors_1_6/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.98f
C928 cp1_buffer_5stage_0/cp1_buffer1_0/charge_pump1_0/capacitors_1_6/capacitor_8_0/capacitor_7_0/buffer_digital_0/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.61f
C929 cp1_buffer_5stage_0/cp1_buffer1_0/charge_pump1_0/capacitors_1_5/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.34f
C930 cp1_buffer_5stage_0/cp1_buffer1_0/charge_pump1_0/capacitors_1_5/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.98f
C931 cp1_buffer_5stage_0/cp1_buffer1_0/charge_pump1_0/capacitors_1_5/capacitor_8_0/capacitor_7_0/buffer_digital_0/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.61f
C932 cp1_buffer_5stage_0/cp1_buffer1_0/charge_pump1_0/capacitors_1_4/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.34f
C933 cp1_buffer_5stage_0/cp1_buffer1_0/charge_pump1_0/capacitors_1_4/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.98f
C934 cp1_buffer_5stage_0/cp1_buffer1_0/charge_pump1_0/capacitors_1_4/capacitor_8_0/capacitor_7_0/buffer_digital_0/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.61f
C935 cp1_buffer_5stage_0/cp1_buffer1_0/charge_pump1_0/capacitors_1_3/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.34f
C936 cp1_buffer_5stage_0/cp1_buffer1_0/charge_pump1_0/capacitors_1_3/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.98f
C937 cp1_buffer_5stage_0/cp1_buffer1_0/charge_pump1_0/capacitors_1_3/capacitor_8_0/capacitor_7_0/buffer_digital_0/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.61f
C938 cp1_buffer_5stage_0/cp1_buffer1_0/charge_pump1_0/capacitors_1_2/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.34f
C939 cp1_buffer_5stage_0/cp1_buffer1_0/charge_pump1_0/capacitors_1_2/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.98f
C940 cp1_buffer_5stage_0/cp1_buffer1_0/charge_pump1_0/capacitors_1_2/capacitor_8_0/capacitor_7_0/buffer_digital_0/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.61f
C941 cp1_buffer_5stage_0/cp1_buffer1_0/charge_pump1_0/capacitors_1_1/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.34f
C942 cp1_buffer_5stage_0/cp1_buffer1_0/charge_pump1_0/capacitors_1_1/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.98f
C943 cp1_buffer_5stage_0/cp1_buffer1_0/charge_pump1_0/capacitors_1_1/capacitor_8_0/capacitor_7_0/buffer_digital_0/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.61f
C944 cp1_buffer_5stage_0/cp1_buffer1_0/charge_pump1_0/capacitors_1_0/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.34f
C945 cp1_buffer_5stage_0/cp1_buffer1_0/charge_pump1_0/capacitors_1_0/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.98f
C946 cp1_buffer_5stage_0/cp1_buffer1_0/charge_pump1_0/capacitors_1_0/capacitor_8_0/capacitor_7_0/buffer_digital_0/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.61f
C947 cp1_buffer_5stage_0/cp1_buffer1_0/charge_pump1_0/capacitor_8_1/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.34f
C948 cp1_buffer_5stage_0/cp1_buffer1_0/charge_pump1_0/clkb cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 89.9f
C949 cp1_buffer_5stage_0/cp1_buffer1_0/charge_pump1_0/capacitor_8_1/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.98f
C950 cp1_buffer_5stage_0/cp1_buffer1_0/charge_pump1_0/capacitor_8_1/capacitor_7_0/buffer_digital_0/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.61f
C951 cp1_buffer_5stage_0/cp1_buffer1_0/charge_pump1_0/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.34f
C952 cp1_buffer_5stage_0/cp1_buffer1_0/charge_pump1_0/clk cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 89f
C953 cp1_buffer_5stage_0/cp1_buffer1_0/charge_pump1_0/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 9.98f
C954 cp1_buffer_5stage_0/cp1_buffer1_0/charge_pump1_0/capacitor_8_0/capacitor_7_0/buffer_digital_0/in cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.61f
C955 cp1_buffer_5stage_0/cp1_buffer1_0/charge_pump1_0/clock_0/a_2432_n962# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 8.68f **FLOATING
C956 cp1_buffer_5stage_0/cp1_buffer1_0/charge_pump1_0/clock_0/a_2020_n482# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.57f **FLOATING
C957 cp1_buffer_5stage_0/cp1_buffer1_0/charge_pump1_0/clock_0/a_344_102# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.81f
C958 cp1_buffer_5stage_0/cp1_buffer1_0/charge_pump1_0/clock_0/a_2402_572# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.17f
C959 cp1_buffer_5stage_0/cp1_buffer1_0/charge_pump1_0/clock_0/a_344_n986# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.38f
C960 cp1_buffer_5stage_0/cp1_buffer1_0/charge_pump1_0/clock_0/a_3246_118# cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 6.83f
C961 cp1_buffer_5stage_0/cp1_buffer1_0/charge_pump1_0/g2 cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.34f
C962 cp1_buffer_5stage_0/cp1_buffer1_0/charge_pump1_0/vin cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 10.4f
C963 scanchain_0/net2 cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.35f
C964 scanchain_0/clkbuf_0_clk/A cp2_buffer_5stage_1/cp2_buffer1_2/charge_pump_0/nmos_diode2_0/VSUBS 2.59f
.ends

