magic
tech sky130A
magscale 1 2
timestamp 1698753667
<< nwell >>
rect -444 1286 460 1468
rect -10 1012 216 1286
rect 1652 -116 1668 0
rect 1652 -318 2756 -116
rect 1654 -320 2756 -318
rect 3928 -320 5062 -34
rect 6570 -164 6584 -6
rect 5484 -346 6584 -164
<< nsubdiff >>
rect 2610 -204 2720 -180
rect 2610 -238 2634 -204
rect 2696 -238 2720 -204
rect 2610 -268 2720 -238
rect 4900 -204 5010 -178
rect 4900 -242 4924 -204
rect 4990 -242 5010 -204
rect 4900 -270 5010 -242
rect 6442 -234 6546 -210
rect 6442 -286 6472 -234
rect 6520 -286 6546 -234
rect 6442 -310 6546 -286
<< nsubdiffcont >>
rect 2634 -238 2696 -204
rect 4924 -242 4990 -204
rect 6472 -286 6520 -234
<< poly >>
rect 692 -32 722 14
rect 884 -32 914 28
rect 1076 -32 1106 30
rect 1268 -32 1298 28
rect 1460 -32 1490 18
rect 1662 2 2746 278
rect 3926 6 4938 106
rect 540 -112 1600 -32
rect 1758 -34 1788 2
rect 1950 -28 1980 2
rect 2142 -28 2172 2
rect 2334 -32 2364 2
rect 2526 -32 2556 2
rect 2996 -38 3026 -4
rect 3188 -38 3218 6
rect 3380 -38 3410 -2
rect 3572 -38 3602 -6
rect 3764 -38 3794 4
rect 4024 -24 4054 6
rect 4216 -30 4246 6
rect 4408 -24 4438 6
rect 4600 -26 4630 6
rect 4792 -24 4822 6
rect 5554 -12 6622 72
rect 540 -178 1598 -112
rect 2848 -266 3800 -38
rect 5586 -46 5616 -12
rect 5778 -46 5808 -12
rect 5970 -40 6000 -12
rect 6162 -40 6192 -12
rect 6354 -50 6384 -12
rect 6842 -38 6872 2
rect 7034 -38 7064 -8
rect 7226 -38 7256 0
rect 7418 -38 7448 4
rect 6656 -300 7498 -38
<< locali >>
rect 1662 252 2746 278
rect 1662 40 1706 252
rect 2658 40 2746 252
rect 1662 2 2746 40
rect 3926 52 4014 106
rect 5554 172 6620 204
rect 4876 52 4938 106
rect 3926 6 4938 52
rect 5554 48 5676 172
rect 6488 48 6620 172
rect 5554 -12 6620 48
rect 540 -66 1598 -38
rect 540 -160 568 -66
rect 1562 -160 1598 -66
rect 540 -178 1598 -160
rect 2848 -80 3800 -50
rect 2610 -204 2720 -180
rect 2610 -240 2634 -204
rect 2696 -240 2720 -204
rect 2610 -268 2720 -240
rect 2848 -246 2886 -80
rect 3778 -246 3800 -80
rect 6656 -108 7498 -46
rect 2848 -266 3800 -246
rect 4900 -204 5008 -176
rect 4900 -242 4924 -204
rect 4990 -242 5008 -204
rect 4900 -270 5008 -242
rect 6442 -234 6546 -210
rect 6442 -286 6472 -234
rect 6520 -286 6546 -234
rect 6442 -310 6546 -286
rect 6656 -242 6672 -108
rect 7456 -242 7498 -108
rect 6656 -300 7498 -242
<< viali >>
rect 1706 40 2658 252
rect 4014 52 4876 320
rect 5676 48 6488 172
rect 568 -160 1562 -66
rect 2634 -238 2696 -204
rect 2634 -240 2696 -238
rect 2886 -246 3778 -80
rect 4924 -242 4990 -204
rect 6472 -286 6520 -234
rect 6672 -242 7456 -108
<< metal1 >>
rect -466 2004 140 2046
rect -466 1532 -418 2004
rect 78 1532 140 2004
rect 2536 1760 3626 1798
rect -466 1366 140 1532
rect -2 996 248 1002
rect -636 948 -518 988
rect -2 942 20 996
rect 238 992 248 996
rect 238 948 262 992
rect 238 942 248 948
rect 0 936 248 942
rect 7200 930 7828 948
rect 7200 870 7216 930
rect 7108 850 7216 870
rect 7608 870 7828 930
rect 7608 850 7938 870
rect 7108 838 7938 850
rect -386 788 -352 836
rect -168 792 -134 836
rect -168 788 -132 792
rect -386 732 -132 788
rect -498 520 108 732
rect -498 48 -446 520
rect 50 48 108 520
rect -498 34 108 48
rect 530 92 1596 534
rect 1662 252 2746 526
rect 530 -2 1600 92
rect 1662 40 1706 252
rect 2658 40 2746 252
rect 1662 2 2746 40
rect 2838 -8 3866 544
rect 3926 320 4946 518
rect 3926 52 4014 320
rect 4876 52 4946 320
rect 3926 6 4946 52
rect 5554 172 6624 542
rect 5554 48 5676 172
rect 6488 48 6624 172
rect 5554 -12 6624 48
rect 6662 0 7498 536
rect 540 -66 1598 -38
rect 540 -160 568 -66
rect 1562 -114 1598 -66
rect 1562 -160 1600 -114
rect 1658 -154 2756 -52
rect 2848 -80 3794 -50
rect 2848 -154 2886 -80
rect 540 -178 1600 -160
rect 568 -256 1600 -178
rect 1640 -204 2886 -154
rect 1640 -240 2634 -204
rect 2696 -240 2886 -204
rect 1640 -246 2886 -240
rect 3778 -154 3794 -80
rect 3926 -154 5062 -36
rect 3778 -204 5062 -154
rect 3778 -242 4924 -204
rect 4990 -242 5062 -204
rect 3778 -246 5062 -242
rect 1640 -304 5062 -246
rect 5478 -234 6548 -52
rect 5478 -286 6472 -234
rect 6520 -286 6548 -234
rect 5478 -290 6548 -286
rect 3926 -322 5062 -304
rect 5484 -336 6548 -290
rect 6656 -108 7498 -38
rect 6656 -242 6672 -108
rect 7456 -242 7498 -108
rect 6656 -300 7498 -242
<< via1 >>
rect -418 1532 78 2004
rect 20 942 238 996
rect 7216 850 7608 930
rect -446 48 50 520
<< metal2 >>
rect -466 2004 140 2046
rect -466 1532 -418 2004
rect 78 1532 140 2004
rect -466 1474 140 1532
rect -660 1070 8996 1082
rect -660 1034 8998 1070
rect -660 928 -612 1034
rect 7406 1030 8998 1034
rect 2 996 248 1002
rect 2 942 20 996
rect 238 992 248 996
rect 238 948 262 992
rect 238 942 248 948
rect 2 936 248 942
rect 7200 930 7634 948
rect 7200 850 7216 930
rect 7608 850 7634 930
rect 7200 838 7634 850
rect -498 520 108 568
rect -498 48 -446 520
rect 50 48 108 520
rect -498 34 108 48
<< via2 >>
rect -418 1532 78 2004
rect 7216 850 7608 930
rect -446 48 50 520
<< metal3 >>
rect -466 2004 140 2046
rect -466 1532 -418 2004
rect 78 1532 140 2004
rect -466 1474 140 1532
rect 7772 1396 8834 1430
rect 7200 930 7634 948
rect -778 798 8 894
rect 7200 850 7216 930
rect 7608 850 7634 930
rect 7200 838 7634 850
rect 7768 946 8834 1396
rect 7768 734 8990 946
rect -498 520 108 568
rect -498 48 -446 520
rect 50 48 108 520
rect 7768 402 8834 734
rect 7772 370 8834 402
rect -498 34 108 48
<< via3 >>
rect -418 1532 78 2004
rect 7216 850 7608 930
rect -446 48 50 520
<< mimcap >>
rect 7800 932 8800 1396
rect 7800 762 7838 932
rect 8118 762 8800 932
rect 7800 402 8800 762
<< mimcapcontact >>
rect 7838 762 8118 932
<< metal4 >>
rect -1378 2004 140 2046
rect -1378 1532 -418 2004
rect 78 1532 140 2004
rect -1378 1474 140 1532
rect -1378 -154 -806 1474
rect 7756 950 8144 954
rect 7200 932 8144 950
rect 7200 930 7838 932
rect 7200 850 7216 930
rect 7608 850 7838 930
rect 7200 838 7838 850
rect 7756 762 7838 838
rect 8118 762 8144 932
rect 7756 726 8144 762
rect -498 520 108 568
rect -498 48 -446 520
rect 50 48 108 520
rect -498 34 108 48
<< via4 >>
rect -446 48 50 520
<< metal5 >>
rect -498 566 108 568
rect -1972 520 108 566
rect -1972 48 -446 520
rect 50 48 108 520
rect -1972 -4 108 48
rect -1972 -6 -60 -4
rect -1972 -154 -1400 -6
use buffer_and_gate  buffer_and_gate_0
timestamp 1698476459
transform 1 0 84 0 1 30
box -116 -30 7470 2020
use buffer_digital  buffer_digital_1 ~/Desktop/charge_pumps2/layout_files
timestamp 1698753667
transform 1 0 -384 0 1 799
box -274 0 415 576
use sky130_fd_pr__nfet_01v8_D4CMYK  sky130_fd_pr__nfet_01v8_D4CMYK_0
timestamp 1698652801
transform 1 0 7097 0 1 40
box -413 -130 413 130
use sky130_fd_pr__nfet_01v8_NJGC45  sky130_fd_pr__nfet_01v8_NJGC45_0
timestamp 1698666719
transform 1 0 1043 0 1 48
box -509 -130 509 130
use sky130_fd_pr__nfet_01v8_NJGC45  sky130_fd_pr__nfet_01v8_NJGC45_1
timestamp 1698666719
transform 1 0 3347 0 1 40
box -509 -130 509 130
use sky130_fd_pr__pfet_01v8_4ZKXAA  sky130_fd_pr__pfet_01v8_4ZKXAA_1
timestamp 1698666719
transform 1 0 4471 0 1 -82
box -545 -142 545 142
use sky130_fd_pr__pfet_01v8_4ZKXAA  sky130_fd_pr__pfet_01v8_4ZKXAA_2
timestamp 1698666719
transform 1 0 6033 0 1 -100
box -545 -142 545 142
use sky130_fd_pr__pfet_01v8_4ZKXAA  sky130_fd_pr__pfet_01v8_4ZKXAA_3
timestamp 1698666719
transform 1 0 2205 0 1 -84
box -545 -142 545 142
<< end >>
