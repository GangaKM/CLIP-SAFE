magic
tech sky130A
magscale 1 2
timestamp 1698914652
<< nwell >>
rect -3654 2366 -2708 2420
rect -3654 1456 -2696 2366
rect -3654 568 -2708 1456
rect -3312 542 -3024 568
rect -3018 556 -2720 568
rect -396 566 184 2640
rect -1728 302 -1042 488
rect -2748 12 -1042 302
rect -1728 10 -1042 12
<< pwell >>
rect -3176 3480 -3114 4296
<< psubdiff >>
rect 426 3536 564 3564
rect 426 3468 460 3536
rect 524 3468 564 3536
rect 426 3440 564 3468
<< nsubdiff >>
rect -18 2512 104 2540
rect -18 2466 10 2512
rect 72 2466 104 2512
rect -18 2430 104 2466
rect -3618 1312 -3498 1338
rect -3618 1250 -3594 1312
rect -3528 1250 -3498 1312
rect -3618 1226 -3498 1250
rect -1502 404 -1394 430
rect -1502 360 -1480 404
rect -1428 360 -1394 404
rect -1502 332 -1394 360
<< psubdiffcont >>
rect 460 3468 524 3536
<< nsubdiffcont >>
rect 10 2466 72 2512
rect -3594 1250 -3528 1312
rect -1480 360 -1428 404
<< poly >>
rect 920 3008 950 3036
rect 822 2970 950 3008
rect 316 2573 449 2603
rect 316 2536 346 2573
rect 2933 2400 2998 2430
rect 2933 2297 2963 2400
rect 3430 2318 3505 2348
rect 3475 2217 3505 2318
rect -3274 1246 -3244 1346
rect -3274 1216 -3208 1246
rect -2800 944 -2720 946
rect -2800 916 -2716 944
rect -2752 816 -2716 916
rect -362 692 -330 790
rect -362 662 -300 692
<< locali >>
rect 444 3536 560 3558
rect 444 3468 458 3536
rect 524 3468 560 3536
rect 444 3448 560 3468
rect -3876 3350 -3688 3430
rect -4052 3322 -2894 3350
rect -4052 3264 -2836 3322
rect -4052 3262 -2894 3264
rect -2908 2916 -2766 2998
rect -2524 2918 -2382 3000
rect 2784 2950 2882 3048
rect 2784 2612 2800 2950
rect 2850 2612 2882 2950
rect -18 2512 104 2540
rect 2784 2520 2882 2612
rect -18 2466 10 2512
rect 72 2466 104 2512
rect -18 2430 104 2466
rect -3618 1312 -3498 1338
rect -3618 1250 -3594 1312
rect -3528 1250 -3498 1312
rect -3618 1226 -3498 1250
rect -1502 404 -1394 430
rect -1502 360 -1480 404
rect -1428 360 -1394 404
rect -1502 332 -1394 360
<< viali >>
rect -3802 4536 4658 4752
rect 458 3468 460 3536
rect 460 3468 524 3536
rect -1684 2750 782 2796
rect 2800 2612 2850 2950
rect 10 2466 72 2512
rect -3594 1250 -3528 1312
rect -1478 360 -1428 404
rect -3800 -654 4732 -378
<< metal1 >>
rect -3835 4752 4779 4979
rect -3835 4536 -3802 4752
rect 4658 4536 4779 4752
rect -3835 4427 4779 4536
rect -3410 4404 640 4427
rect -4134 3600 -3658 3612
rect -4134 3570 -3548 3600
rect -3862 3540 -3548 3570
rect -3862 3536 -3630 3540
rect -3640 3458 -3630 3536
rect -3558 3458 -3548 3540
rect -3410 2770 -3346 4404
rect -3264 4326 -3224 4404
rect -3266 3706 -3224 4326
rect -3266 3702 -3226 3706
rect -3186 3554 -3176 4370
rect -3114 3554 -3104 4370
rect -3068 4323 -3028 4404
rect -3068 3608 -3024 4323
rect 312 4312 640 4404
rect 452 3536 530 3548
rect 38 3452 48 3506
rect 152 3452 162 3506
rect 452 3468 458 3536
rect 524 3468 530 3536
rect 452 3456 530 3468
rect 458 3408 524 3456
rect 3588 3442 3598 3500
rect 3704 3442 3714 3500
rect 3867 3470 4507 3507
rect -946 3160 -936 3216
rect -754 3186 -744 3216
rect -754 3160 -672 3186
rect -780 3112 -672 3160
rect -203 3139 -114 3149
rect -786 3084 -680 3096
rect -786 3068 -682 3084
rect -210 3052 -200 3139
rect -134 3052 -114 3139
rect 6 3114 36 3340
rect 232 3258 712 3408
rect 382 3246 680 3258
rect 132 3156 958 3204
rect 2 3054 998 3114
rect -203 3042 -114 3052
rect 1119 3046 1218 3048
rect -1466 2972 -1456 3028
rect -1274 2972 -1264 3028
rect 50 2968 876 3016
rect 1086 2986 1218 3046
rect 810 2932 852 2968
rect 1086 2932 1181 2986
rect -14 2872 1181 2932
rect 1119 2871 1181 2872
rect 2784 2950 2882 3048
rect 2976 3042 2986 3149
rect 3075 3042 3085 3149
rect -1684 2802 794 2822
rect -3410 2690 -3300 2770
rect -1696 2750 -1684 2802
rect 784 2750 794 2802
rect -1696 2744 794 2750
rect -1696 2730 772 2744
rect -3606 1312 -3516 1318
rect -3410 1312 -3346 2690
rect -2630 2689 -1692 2702
rect -2755 2572 -2702 2679
rect -2640 2629 -2630 2689
rect -2002 2629 -1692 2689
rect 523 2653 1227 2699
rect 1702 2653 1887 2699
rect -650 2542 -556 2590
rect -362 2530 -330 2592
rect -2 2570 1038 2622
rect -2 2568 90 2570
rect -3296 2246 -3256 2328
rect -3296 2194 -3252 2246
rect -3606 1250 -3594 1312
rect -3528 1250 -3346 1312
rect -3292 1618 -3252 2194
rect -3292 1348 -3264 1618
rect -3292 1304 -3244 1348
rect -3606 1244 -3516 1250
rect -3410 496 -3346 1250
rect -3284 720 -3244 1304
rect -3182 730 -3124 2292
rect -3074 2142 -2934 2344
rect -3084 1514 -2934 2142
rect -3194 584 -3124 730
rect -3074 634 -2934 1514
rect -3072 622 -3032 634
rect -3194 496 -3128 584
rect -2870 496 -2812 2344
rect -366 2302 -328 2530
rect -479 2249 -406 2299
rect -372 2244 -322 2302
rect -2760 2202 -2708 2210
rect -2768 796 -2758 2202
rect -2694 796 -2684 2202
rect -372 2138 -321 2244
rect -371 2083 -321 2138
rect -270 2148 -212 2566
rect -204 2534 90 2568
rect -22 2520 90 2534
rect 834 2522 1070 2524
rect -22 2512 108 2520
rect -22 2466 10 2512
rect 72 2468 108 2512
rect 186 2468 1070 2522
rect 72 2466 84 2468
rect -22 2462 84 2466
rect -2 2460 84 2462
rect 186 2458 292 2468
rect 834 2466 1070 2468
rect 1181 2473 1227 2653
rect 1841 2614 1887 2653
rect 2784 2612 2800 2950
rect 2868 2612 2882 2950
rect 2784 2520 2882 2612
rect 186 2450 264 2458
rect -152 2410 -112 2434
rect -158 2380 -102 2410
rect -152 2324 -112 2380
rect -160 2250 -110 2324
rect 186 2250 234 2450
rect 1181 2427 1869 2473
rect 298 2410 936 2422
rect 280 2380 936 2410
rect 298 2370 936 2380
rect 1823 2378 1869 2427
rect 1804 2326 1910 2378
rect 2150 2334 2160 2408
rect 2266 2334 2276 2408
rect 2918 2278 2966 2734
rect -160 2202 234 2250
rect -476 1508 -400 1556
rect -366 750 -324 2083
rect -270 2010 -216 2148
rect -160 2028 -110 2202
rect 3008 2194 3066 2768
rect 3112 2346 3156 2654
rect 3268 2346 3304 2734
rect 3112 2310 3306 2346
rect 3112 2198 3156 2310
rect -366 746 -328 750
rect -270 612 -206 2010
rect -152 700 -112 2028
rect -152 656 54 700
rect -260 496 -206 612
rect -3924 404 -112 496
rect -3924 360 -1478 404
rect -1428 360 -112 404
rect -3924 346 -112 360
rect -3924 340 -2354 346
rect -1338 340 -112 346
rect -3412 295 -3344 340
rect -3845 257 -2947 295
rect -2803 294 -2371 295
rect -3845 84 -3807 257
rect -3590 240 -2948 257
rect -2803 246 -1128 294
rect -2803 245 -2371 246
rect -3728 130 -2922 194
rect -3690 84 -3048 94
rect -3845 46 -3048 84
rect -3690 44 -3048 46
rect -2964 -256 -2926 130
rect -2803 104 -2753 245
rect -1100 192 -1062 340
rect -1028 338 -112 340
rect -724 273 -676 338
rect -1130 186 -1062 192
rect -2694 130 -1062 186
rect -975 223 -107 273
rect -2694 126 -1066 130
rect -2806 66 -2753 104
rect -975 72 -925 223
rect -94 176 -56 190
rect -872 126 -52 176
rect -2666 66 -1342 70
rect -2806 22 -1342 66
rect -975 22 -186 72
rect -2806 16 -2624 22
rect -2806 -256 -2754 16
rect -1420 -256 -1382 -254
rect -94 -256 -56 126
rect 10 -256 54 656
rect 1818 -256 2110 2060
rect 3008 2022 3068 2194
rect 3348 2026 3412 2782
rect 3536 2634 3569 3060
rect 3462 2598 3569 2634
rect 3462 2218 3498 2598
rect 3536 2178 3569 2598
rect -3834 -372 4728 -256
rect -3834 -378 4744 -372
rect -3834 -654 -3800 -378
rect 4732 -654 4744 -378
rect -3834 -660 4744 -654
rect -3834 -770 4728 -660
<< via1 >>
rect -3802 4536 4658 4752
rect -3630 3458 -3558 3540
rect -3176 3554 -3114 4370
rect 48 3452 152 3506
rect 3598 3442 3704 3500
rect -936 3160 -754 3216
rect -200 3052 -134 3139
rect -1456 2972 -1274 3028
rect 2986 3042 3075 3149
rect -1684 2796 784 2802
rect -1684 2750 782 2796
rect 782 2750 784 2796
rect -2630 2629 -2002 2689
rect -2758 796 -2694 2202
rect 2800 2612 2850 2950
rect 2850 2612 2868 2950
rect 2160 2334 2266 2408
rect -3800 -654 4732 -378
<< metal2 >>
rect -3835 4752 4779 4979
rect -3835 4536 -3802 4752
rect 4658 4536 4779 4752
rect -3835 4427 4779 4536
rect -3176 4370 -3114 4380
rect -3630 3540 -3558 3550
rect -3630 3448 -3558 3458
rect -3176 3423 -3114 3554
rect 48 3506 152 3516
rect 48 3442 52 3452
rect 142 3442 152 3452
rect 3598 3500 3704 3510
rect 52 3430 142 3440
rect 3598 3432 3704 3442
rect -3176 3361 -2815 3423
rect -936 3216 -754 3226
rect -936 3150 -754 3160
rect -203 3151 -114 3161
rect -1456 3028 -1274 3038
rect -203 3034 -114 3044
rect 2986 3149 3075 3159
rect 2986 3032 3075 3042
rect -1456 2962 -1274 2972
rect 2800 2950 2868 2960
rect -1684 2808 784 2818
rect -3564 2750 -1684 2808
rect -3564 2748 784 2750
rect -1684 2740 784 2748
rect -2630 2691 -2002 2699
rect -3583 2689 -2002 2691
rect -3583 2629 -2630 2689
rect -3583 2621 -2002 2629
rect -2630 2619 -2002 2621
rect 2800 2602 2868 2612
rect 1994 2502 2094 2541
rect 2320 2502 2407 2541
rect 2160 2408 2266 2418
rect 2160 2324 2266 2334
rect -2758 2210 -2694 2212
rect -2768 2202 -2694 2210
rect -2768 796 -2758 2202
rect 4256 1738 4712 1826
rect -2768 786 -2694 796
rect -2768 -256 -2698 786
rect -3800 -368 4728 -256
rect -3800 -378 4732 -368
rect -3800 -664 4732 -654
rect -3800 -770 4728 -664
<< via2 >>
rect -3802 4536 4658 4752
rect -3630 3458 -3558 3540
rect 52 3452 142 3506
rect 52 3440 142 3452
rect 3598 3442 3704 3500
rect -936 3160 -754 3216
rect -203 3139 -114 3151
rect -203 3052 -200 3139
rect -200 3052 -134 3139
rect -134 3052 -114 3139
rect -203 3044 -114 3052
rect 2986 3042 3075 3149
rect -1456 2972 -1274 3028
rect -1684 2802 784 2808
rect -1684 2750 784 2802
rect 2800 2612 2868 2950
rect 2160 2334 2266 2408
<< metal3 >>
rect -3835 4766 4779 4979
rect -3835 4494 -3802 4766
rect 4654 4752 4779 4766
rect 4658 4536 4779 4752
rect 4654 4494 4779 4536
rect -3835 4427 4779 4494
rect -3640 3540 -3548 3545
rect -3640 3458 -3630 3540
rect -3558 3530 -3548 3540
rect -3558 3464 -138 3530
rect -3558 3458 -3548 3464
rect -3640 3453 -3548 3458
rect -960 3223 -780 3224
rect -3569 3216 -743 3223
rect -3569 3160 -936 3216
rect -754 3160 -743 3216
rect -3569 3154 -743 3160
rect -204 3156 -138 3464
rect 32 3506 166 3512
rect 32 3440 52 3506
rect 142 3440 166 3506
rect 32 3434 166 3440
rect 386 3500 3715 3508
rect 386 3442 3598 3500
rect 3704 3442 3715 3500
rect 386 3434 3715 3442
rect -213 3155 -104 3156
rect -213 3151 -26 3155
rect -213 3044 -203 3151
rect -114 3138 -26 3151
rect 2976 3149 3085 3154
rect 2976 3138 2986 3149
rect -114 3050 2986 3138
rect -114 3044 -26 3050
rect -213 3040 -26 3044
rect 2976 3042 2986 3050
rect 3075 3042 3085 3149
rect -213 3039 -104 3040
rect 2976 3037 3085 3042
rect -1466 3028 -1264 3033
rect -1466 3024 -1456 3028
rect -3558 2972 -1456 3024
rect -1274 2972 -1264 3028
rect -3558 2967 -1264 2972
rect -3558 2961 -1330 2967
rect -1510 2956 -1330 2961
rect 2790 2950 2878 2955
rect -1684 2813 794 2822
rect -1694 2808 794 2813
rect -1694 2800 -1684 2808
rect -1726 2750 -1684 2800
rect 784 2750 794 2808
rect -1726 2745 794 2750
rect -1726 2732 768 2745
rect 700 2534 768 2732
rect 2790 2612 2800 2950
rect 2868 2698 2878 2950
rect 4301 2698 4387 4427
rect 2868 2612 4387 2698
rect 2790 2607 2878 2612
rect 700 2466 2270 2534
rect 2150 2413 2270 2466
rect 2150 2408 2276 2413
rect 2150 2334 2160 2408
rect 2266 2334 2276 2408
rect 2150 2329 2276 2334
rect 2202 2322 2270 2329
rect 809 2196 4482 2257
rect 809 2182 1764 2196
rect 2138 2182 4482 2196
<< via3 >>
rect -3802 4752 4654 4766
rect -3802 4536 4658 4752
rect -3802 4494 4654 4536
<< metal4 >>
rect -3835 4766 4779 4979
rect -3835 4494 -3802 4766
rect 4654 4752 4779 4766
rect 4658 4536 4779 4752
rect 4654 4494 4779 4536
rect -3835 4427 4779 4494
use firststage_compact  firststage_compact_0
timestamp 1698871213
transform 1 0 -43 0 1 -468
box -3293 1004 775 4931
use integrator_full_new_compact  integrator_full_new_compact_0
timestamp 1698861754
transform 1 0 386 0 1 3329
box -386 -3496 4003 1133
use sky130_fd_pr__nfet_01v8_5WVHMA  sky130_fd_pr__nfet_01v8_5WVHMA_0
timestamp 1698873245
transform 0 -1 3040 1 0 2463
box -317 -130 317 130
use sky130_fd_pr__nfet_01v8_5WVHMA  sky130_fd_pr__nfet_01v8_5WVHMA_1
timestamp 1698873245
transform 0 -1 3384 1 0 2477
box -317 -130 317 130
use sky130_fd_pr__nfet_01v8_53744R  sky130_fd_pr__nfet_01v8_53744R_0
timestamp 1698787694
transform 0 -1 -3778 1 0 3494
box -246 -310 246 310
use sky130_fd_pr__nfet_01v8_FU3CJE  sky130_fd_pr__nfet_01v8_FU3CJE_0
timestamp 1698611618
transform 1 0 503 0 1 3086
box -509 -130 509 130
use sky130_fd_pr__nfet_01v8_GWAZJ9  sky130_fd_pr__nfet_01v8_GWAZJ9_0
timestamp 1698873245
transform 1 0 -3323 0 1 164
box -413 -130 413 130
use sky130_fd_pr__nfet_01v8_GWAZJ9  sky130_fd_pr__nfet_01v8_GWAZJ9_1
timestamp 1698873245
transform 1 0 -469 0 1 152
box -413 -130 413 130
use sky130_fd_pr__nfet_01v8_GWAZJ9  sky130_fd_pr__nfet_01v8_GWAZJ9_2
timestamp 1698873245
transform 1 0 667 0 1 2494
box -413 -130 413 130
use sky130_fd_pr__nfet_01v8_GWXQMW  sky130_fd_pr__nfet_01v8_GWXQMW_0
timestamp 1698611618
transform 0 -1 -3146 1 0 3969
box -413 -130 413 130
use sky130_fd_pr__pfet_01v8_ACB9FB  sky130_fd_pr__pfet_01v8_ACB9FB_0
timestamp 1698611618
transform 0 -1 -3156 1 0 991
box -449 -142 449 142
use sky130_fd_pr__pfet_01v8_ACB9FB  sky130_fd_pr__pfet_01v8_ACB9FB_1
timestamp 1698611618
transform 0 -1 -3166 1 0 1883
box -449 -142 449 142
use sky130_fd_pr__pfet_01v8_ACB9FB  sky130_fd_pr__pfet_01v8_ACB9FB_2
timestamp 1698611618
transform 0 -1 -2840 1 0 1171
box -449 -142 449 142
use sky130_fd_pr__pfet_01v8_ACB9FB  sky130_fd_pr__pfet_01v8_ACB9FB_3
timestamp 1698611618
transform 0 -1 -2840 1 0 1939
box -449 -142 449 142
use sky130_fd_pr__pfet_01v8_DCBZKP  sky130_fd_pr__pfet_01v8_DCBZKP_0
timestamp 1698611618
transform 1 0 -1896 0 1 158
box -848 -142 848 142
use sky130_fd_pr__pfet_01v8_WMSBVE  sky130_fd_pr__pfet_01v8_WMSBVE_0
timestamp 1698611618
transform 0 -1 -240 1 0 1589
box -1025 -142 1025 142
<< labels >>
rlabel metal4 -3652 4448 -3652 4448 1 Vdd
rlabel metal1 -598 2574 -598 2574 1 Vbp
rlabel metal3 3108 3462 3108 3462 1 Vcmref
rlabel metal3 -3509 3189 -3509 3189 1 Vbias
rlabel metal3 -3509 2980 -3509 2980 1 Vs
rlabel metal2 -3490 2771 -3490 2771 1 vd2
rlabel metal2 -3506 2656 -3506 2656 1 vd1
rlabel metal1 4425 3485 4425 3485 1 Vcmref
rlabel metal2 4641 1770 4641 1770 1 vo1
rlabel space 4480 2009 6100 2501 1 ete
rlabel metal1 -4110 3584 -4110 3584 1 Vbias_int
<< end >>
