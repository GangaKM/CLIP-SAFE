magic
tech sky130A
magscale 1 2
timestamp 1698837886
<< nwell >>
rect -449 104 545 142
rect -545 -104 545 104
rect -545 -142 449 -104
<< pmos >>
rect -447 -42 -417 42
rect -351 -42 -321 42
rect -255 -42 -225 42
rect -159 -42 -129 42
rect -63 -42 -33 42
rect 33 -42 63 42
rect 129 -42 159 42
rect 225 -42 255 42
rect 321 -42 351 42
rect 417 -42 447 42
<< pdiff >>
rect -509 30 -447 42
rect -509 -30 -497 30
rect -463 -30 -447 30
rect -509 -42 -447 -30
rect -417 30 -351 42
rect -417 -30 -401 30
rect -367 -30 -351 30
rect -417 -42 -351 -30
rect -321 30 -255 42
rect -321 -30 -305 30
rect -271 -30 -255 30
rect -321 -42 -255 -30
rect -225 30 -159 42
rect -225 -30 -209 30
rect -175 -30 -159 30
rect -225 -42 -159 -30
rect -129 30 -63 42
rect -129 -30 -113 30
rect -79 -30 -63 30
rect -129 -42 -63 -30
rect -33 30 33 42
rect -33 -30 -17 30
rect 17 -30 33 30
rect -33 -42 33 -30
rect 63 30 129 42
rect 63 -30 79 30
rect 113 -30 129 30
rect 63 -42 129 -30
rect 159 30 225 42
rect 159 -30 175 30
rect 209 -30 225 30
rect 159 -42 225 -30
rect 255 30 321 42
rect 255 -30 271 30
rect 305 -30 321 30
rect 255 -42 321 -30
rect 351 30 417 42
rect 351 -30 367 30
rect 401 -30 417 30
rect 351 -42 417 -30
rect 447 30 509 42
rect 447 -30 463 30
rect 497 -30 509 30
rect 447 -42 509 -30
<< pdiffc >>
rect -497 -30 -463 30
rect -401 -30 -367 30
rect -305 -30 -271 30
rect -209 -30 -175 30
rect -113 -30 -79 30
rect -17 -30 17 30
rect 79 -30 113 30
rect 175 -30 209 30
rect 271 -30 305 30
rect 367 -30 401 30
rect 463 -30 497 30
<< poly >>
rect -369 123 -303 139
rect -369 89 -353 123
rect -319 89 -303 123
rect -369 73 -303 89
rect -177 123 -111 139
rect -177 89 -161 123
rect -127 89 -111 123
rect -177 73 -111 89
rect 15 123 81 139
rect 15 89 31 123
rect 65 89 81 123
rect 15 73 81 89
rect 207 123 273 139
rect 207 89 223 123
rect 257 89 273 123
rect 207 73 273 89
rect 399 123 465 139
rect 399 89 415 123
rect 449 89 465 123
rect 399 73 465 89
rect -447 42 -417 68
rect -351 42 -321 73
rect -255 42 -225 68
rect -159 42 -129 73
rect -63 42 -33 68
rect 33 42 63 73
rect 129 42 159 68
rect 225 42 255 73
rect 321 42 351 68
rect 417 42 447 73
rect -447 -73 -417 -42
rect -351 -68 -321 -42
rect -255 -73 -225 -42
rect -159 -68 -129 -42
rect -63 -73 -33 -42
rect 33 -68 63 -42
rect 129 -73 159 -42
rect 225 -68 255 -42
rect 321 -73 351 -42
rect 417 -68 447 -42
rect -465 -89 -399 -73
rect -465 -123 -449 -89
rect -415 -123 -399 -89
rect -465 -139 -399 -123
rect -273 -89 -207 -73
rect -273 -123 -257 -89
rect -223 -123 -207 -89
rect -273 -139 -207 -123
rect -81 -89 -15 -73
rect -81 -123 -65 -89
rect -31 -123 -15 -89
rect -81 -139 -15 -123
rect 111 -89 177 -73
rect 111 -123 127 -89
rect 161 -123 177 -89
rect 111 -139 177 -123
rect 303 -89 369 -73
rect 303 -123 319 -89
rect 353 -123 369 -89
rect 303 -139 369 -123
<< polycont >>
rect -353 89 -319 123
rect -161 89 -127 123
rect 31 89 65 123
rect 223 89 257 123
rect 415 89 449 123
rect -449 -123 -415 -89
rect -257 -123 -223 -89
rect -65 -123 -31 -89
rect 127 -123 161 -89
rect 319 -123 353 -89
<< locali >>
rect -369 89 -353 123
rect -319 89 -303 123
rect -177 89 -161 123
rect -127 89 -111 123
rect 15 89 31 123
rect 65 89 81 123
rect 207 89 223 123
rect 257 89 273 123
rect 399 89 415 123
rect 449 89 465 123
rect -497 30 -463 46
rect -497 -46 -463 -30
rect -401 30 -367 46
rect -401 -46 -367 -30
rect -305 30 -271 46
rect -305 -46 -271 -30
rect -209 30 -175 46
rect -209 -46 -175 -30
rect -113 30 -79 46
rect -113 -46 -79 -30
rect -17 30 17 46
rect -17 -46 17 -30
rect 79 30 113 46
rect 79 -46 113 -30
rect 175 30 209 46
rect 175 -46 209 -30
rect 271 30 305 46
rect 271 -46 305 -30
rect 367 30 401 46
rect 367 -46 401 -30
rect 463 30 497 46
rect 463 -46 497 -30
rect -465 -123 -449 -89
rect -415 -123 -399 -89
rect -273 -123 -257 -89
rect -223 -123 -207 -89
rect -81 -123 -65 -89
rect -31 -123 -15 -89
rect 111 -123 127 -89
rect 161 -123 177 -89
rect 303 -123 319 -89
rect 353 -123 369 -89
<< viali >>
rect -497 -30 -463 30
rect -401 -30 -367 30
rect -305 -30 -271 30
rect -209 -30 -175 30
rect -113 -30 -79 30
rect -17 -30 17 30
rect 79 -30 113 30
rect 175 -30 209 30
rect 271 -30 305 30
rect 367 -30 401 30
rect 463 -30 497 30
<< metal1 >>
rect -503 30 -457 42
rect -503 -30 -497 30
rect -463 -30 -457 30
rect -503 -42 -457 -30
rect -407 30 -361 42
rect -407 -30 -401 30
rect -367 -30 -361 30
rect -407 -42 -361 -30
rect -311 30 -265 42
rect -311 -30 -305 30
rect -271 -30 -265 30
rect -311 -42 -265 -30
rect -215 30 -169 42
rect -215 -30 -209 30
rect -175 -30 -169 30
rect -215 -42 -169 -30
rect -119 30 -73 42
rect -119 -30 -113 30
rect -79 -30 -73 30
rect -119 -42 -73 -30
rect -23 30 23 42
rect -23 -30 -17 30
rect 17 -30 23 30
rect -23 -42 23 -30
rect 73 30 119 42
rect 73 -30 79 30
rect 113 -30 119 30
rect 73 -42 119 -30
rect 169 30 215 42
rect 169 -30 175 30
rect 209 -30 215 30
rect 169 -42 215 -30
rect 265 30 311 42
rect 265 -30 271 30
rect 305 -30 311 30
rect 265 -42 311 -30
rect 361 30 407 42
rect 361 -30 367 30
rect 401 -30 407 30
rect 361 -42 407 -30
rect 457 30 503 42
rect 457 -30 463 30
rect 497 -30 503 30
rect 457 -42 503 -30
<< properties >>
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 0.42 l 0.15 m 1 nf 10 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 0 botc 0 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 0 viasrc 100 viadrn 100 viagate 0 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
