magic
tech sky130A
magscale 1 2
timestamp 1698651669
<< psubdiff >>
rect 5661 -409 5748 -383
rect 5661 -450 5688 -409
rect 5722 -450 5748 -409
rect 5661 -475 5748 -450
<< psubdiffcont >>
rect 5688 -450 5722 -409
<< poly >>
rect 38 -356 173 -322
rect 38 -375 72 -356
rect 932 -359 1061 -329
rect 932 -402 962 -359
rect 1890 -362 2013 -332
rect 2848 -352 2977 -322
rect 3830 -329 3860 -324
rect 1890 -394 1920 -362
rect 2848 -384 2878 -352
rect 3830 -359 3959 -329
rect 4772 -356 4901 -326
rect 3830 -386 3860 -359
rect 4772 -388 4802 -356
<< locali >>
rect 302 -290 988 -258
rect 5661 -409 5748 -383
rect 5661 -451 5687 -409
rect 5722 -451 5748 -409
rect 5661 -475 5748 -451
rect -16 -612 5796 -526
rect -16 -614 666 -612
<< viali >>
rect 5687 -450 5688 -409
rect 5688 -450 5722 -409
rect 5687 -451 5722 -450
<< metal1 >>
rect -224 1534 6008 1598
rect -242 1330 -232 1534
rect 5994 1330 6008 1534
rect -224 1244 6008 1330
rect 424 1064 528 1244
rect 5503 1228 5623 1244
rect 5740 1217 5856 1244
rect -274 960 914 1064
rect -274 -578 -170 960
rect 424 930 528 960
rect 870 244 974 258
rect 870 190 882 244
rect 954 190 974 244
rect 1254 192 1264 250
rect 1346 192 1356 250
rect 2424 192 2434 252
rect 2508 192 2518 252
rect 2812 190 2822 248
rect 2892 190 2902 248
rect 870 188 974 190
rect -12 -432 16 -212
rect 302 -290 988 -264
rect 124 -360 740 -326
rect 882 -420 916 -290
rect 1014 -376 1646 -326
rect 1840 -416 1874 -260
rect 1968 -372 2600 -322
rect -14 -460 790 -432
rect -12 -470 16 -460
rect 878 -472 1680 -420
rect 1840 -454 2646 -416
rect 1844 -468 2646 -454
rect 2794 -424 2828 -260
rect 2934 -372 3560 -330
rect 3780 -424 3814 -266
rect 3920 -376 4546 -334
rect 4722 -420 4756 -274
rect 4854 -374 5480 -332
rect 5680 -397 5728 -213
rect 5680 -409 5730 -397
rect 2794 -476 3596 -424
rect 3778 -476 4580 -424
rect 4720 -472 5522 -420
rect 5680 -451 5687 -409
rect 5722 -451 5730 -409
rect 5680 -464 5730 -451
rect 26 -520 664 -516
rect -16 -526 666 -520
rect -16 -578 5796 -526
rect -274 -612 5796 -578
rect -274 -614 666 -612
rect -274 -682 2 -614
rect 826 -1442 836 -1378
rect 926 -1442 936 -1378
rect 1212 -1440 1222 -1376
rect 1312 -1440 1322 -1376
rect 2366 -1386 2480 -1372
rect 2366 -1442 2404 -1386
rect 2472 -1442 2482 -1386
rect 2366 -1444 2480 -1442
rect 2778 -1444 2788 -1390
rect 2852 -1444 2862 -1390
rect -170 -1820 5588 -1818
rect 5864 -1820 5962 -178
rect -170 -1890 6052 -1820
rect -146 -1936 6052 -1890
rect -154 -2114 -144 -1936
rect 6022 -2114 6052 -1936
rect -146 -2214 6052 -2114
<< via1 >>
rect -232 1330 5994 1534
rect 882 190 954 244
rect 1264 192 1346 250
rect 2434 192 2508 252
rect 2822 190 2892 248
rect 836 -1442 926 -1378
rect 1222 -1440 1312 -1376
rect 2404 -1442 2472 -1386
rect 2788 -1444 2852 -1390
rect -144 -2114 6022 -1936
<< metal2 >>
rect -232 1534 5994 1544
rect -232 1320 5994 1330
rect -431 296 1314 326
rect 1284 262 1314 296
rect 870 244 974 258
rect 870 224 882 244
rect -436 190 882 224
rect 954 190 974 244
rect 1258 250 1358 262
rect 1258 192 1264 250
rect 1346 192 1358 250
rect 1258 190 1358 192
rect 2434 252 2508 262
rect -436 188 974 190
rect 882 180 954 188
rect 1264 182 1346 190
rect 2434 182 2508 192
rect 2822 248 2892 258
rect 2822 180 2892 190
rect 4746 -80 4874 -70
rect 4746 -166 4874 -156
rect -300 -1318 1284 -1286
rect 776 -1366 954 -1364
rect 1252 -1366 1284 -1318
rect 776 -1378 956 -1366
rect 776 -1424 836 -1378
rect -308 -1442 836 -1424
rect 926 -1442 956 -1378
rect -308 -1446 956 -1442
rect 1174 -1376 1334 -1366
rect 1174 -1440 1222 -1376
rect 1312 -1440 1334 -1376
rect 1174 -1446 1334 -1440
rect 2366 -1382 2480 -1372
rect 2366 -1442 2404 -1382
rect 2472 -1442 2480 -1382
rect 2366 -1444 2480 -1442
rect 2788 -1384 2852 -1374
rect -308 -1452 954 -1446
rect 1222 -1450 1312 -1446
rect 2404 -1452 2472 -1444
rect 2788 -1454 2852 -1444
rect 4718 -1712 4846 -1702
rect 4718 -1800 4846 -1790
rect -144 -1936 6022 -1926
rect -144 -2124 6022 -2114
<< via2 >>
rect -232 1330 5994 1534
rect 2434 192 2508 252
rect 2822 190 2892 248
rect 4746 -156 4874 -80
rect 2404 -1386 2472 -1382
rect 2404 -1438 2472 -1386
rect 2788 -1390 2852 -1384
rect 2788 -1444 2852 -1390
rect 4718 -1790 4846 -1712
rect -144 -2114 6022 -1936
<< metal3 >>
rect -242 1294 -232 1576
rect 6000 1294 6010 1576
rect -460 388 2506 460
rect 2434 274 2506 388
rect 2410 252 2528 274
rect 2410 192 2434 252
rect 2508 192 2528 252
rect 2410 184 2528 192
rect 2796 248 2914 274
rect 2796 190 2822 248
rect 2892 190 2914 248
rect 2796 184 2914 190
rect 2812 -80 2892 184
rect -435 -128 2892 -80
rect 4736 -80 4884 -75
rect -435 -158 2890 -128
rect 4736 -156 4746 -80
rect 4874 -82 4884 -80
rect 4874 -152 6449 -82
rect 4874 -156 4944 -152
rect 4736 -161 4884 -156
rect -321 -1235 2462 -1173
rect 2400 -1356 2462 -1235
rect 2366 -1382 2482 -1356
rect 2798 -1358 2858 -1356
rect 2366 -1438 2404 -1382
rect 2472 -1438 2482 -1382
rect 2366 -1444 2482 -1438
rect 2772 -1384 2886 -1358
rect 2772 -1444 2788 -1384
rect 2852 -1444 2886 -1384
rect 2772 -1450 2886 -1444
rect 2798 -1732 2858 -1450
rect -320 -1792 2858 -1732
rect 4708 -1712 4856 -1707
rect 4708 -1790 4718 -1712
rect 4846 -1780 6436 -1712
rect 4846 -1790 4856 -1780
rect 4708 -1795 4856 -1790
rect -154 -2114 -144 -1896
rect 6018 -1931 6028 -1896
rect 6018 -1936 6032 -1931
rect 6022 -2114 6032 -1936
rect -154 -2119 6032 -2114
<< via3 >>
rect -232 1534 6000 1576
rect -232 1330 5994 1534
rect 5994 1330 6000 1534
rect -232 1294 6000 1330
rect -144 -1936 6018 -1896
rect -144 -2114 6018 -1936
<< metal4 >>
rect -232 1577 6022 1614
rect -233 1576 6022 1577
rect -233 1294 -232 1576
rect 6000 1294 6022 1576
rect -233 1293 6022 1294
rect -232 1228 6022 1293
rect -232 1214 4944 1228
rect 5714 1214 6022 1228
rect -145 -1896 -128 -1895
rect -145 -2114 -144 -1896
rect -145 -2115 -128 -2114
<< via4 >>
rect -128 -1896 6024 -1892
rect -128 -2114 6018 -1896
rect 6018 -2114 6024 -1896
rect -128 -2174 6024 -2114
<< metal5 >>
rect 5618 -1818 6050 -1814
rect -146 -1868 6050 -1818
rect -152 -1892 6050 -1868
rect -152 -2174 -128 -1892
rect 6024 -2174 6050 -1892
rect -152 -2198 6050 -2174
rect -146 -2214 6050 -2198
use comparator_full_compact  comparator_full_compact_0
timestamp 1698651669
transform 1 0 622 0 1 -292
box -794 -4 5299 1494
use comparator_full_compact  comparator_full_compact_1
timestamp 1698651669
transform 1 0 592 0 1 -1922
box -794 -4 5299 1494
use reference  reference_0
timestamp 1698586885
transform 1 0 -2146 0 1 -1085
box -66 -1120 1956 620
use sky130_fd_pr__nfet_01v8_GWFSUW  sky130_fd_pr__nfet_01v8_GWFSUW_0
timestamp 1698622134
transform 1 0 389 0 1 -442
box -413 -130 413 130
use sky130_fd_pr__nfet_01v8_GWFSUW  sky130_fd_pr__nfet_01v8_GWFSUW_1
timestamp 1698622134
transform 1 0 1283 0 1 -446
box -413 -130 413 130
use sky130_fd_pr__nfet_01v8_GWFSUW  sky130_fd_pr__nfet_01v8_GWFSUW_2
timestamp 1698622134
transform 1 0 2241 0 1 -444
box -413 -130 413 130
use sky130_fd_pr__nfet_01v8_GWFSUW  sky130_fd_pr__nfet_01v8_GWFSUW_3
timestamp 1698622134
transform 1 0 3199 0 1 -444
box -413 -130 413 130
use sky130_fd_pr__nfet_01v8_GWFSUW  sky130_fd_pr__nfet_01v8_GWFSUW_4
timestamp 1698622134
transform 1 0 4181 0 1 -446
box -413 -130 413 130
use sky130_fd_pr__nfet_01v8_GWFSUW  sky130_fd_pr__nfet_01v8_GWFSUW_5
timestamp 1698622134
transform 1 0 5123 0 1 -446
box -413 -130 413 130
<< labels >>
rlabel metal2 -258 -1435 -258 -1435 1 Vc-
rlabel metal2 -253 -1302 -253 -1302 1 V+
rlabel metal3 -289 -1211 -289 -1211 1 V-
rlabel metal3 -298 -1760 -298 -1760 1 Vc+
rlabel metal3 -373 430 -373 430 1 V-
rlabel metal2 -369 312 -369 312 1 V+
rlabel metal2 -380 200 -380 200 1 Vc+
rlabel metal3 -358 -112 -358 -112 1 Vc-
rlabel metal3 6269 -129 6269 -129 1 Q2
rlabel metal3 6329 -1756 6329 -1756 1 Q
<< end >>
