magic
tech sky130A
magscale 1 2
timestamp 1698771642
<< viali >>
rect 6653 8585 6687 8619
rect 1501 8449 1535 8483
rect 3617 8449 3651 8483
rect 6745 8449 6779 8483
rect 7481 8381 7515 8415
rect 1685 8313 1719 8347
rect 6929 8313 6963 8347
rect 2329 8245 2363 8279
rect 5181 8041 5215 8075
rect 5273 7905 5307 7939
rect 1501 7837 1535 7871
rect 2697 7837 2731 7871
rect 2881 7837 2915 7871
rect 4537 7837 4571 7871
rect 4905 7837 4939 7871
rect 7297 7837 7331 7871
rect 4997 7769 5031 7803
rect 5181 7769 5215 7803
rect 5549 7769 5583 7803
rect 1593 7701 1627 7735
rect 2973 7701 3007 7735
rect 4721 7701 4755 7735
rect 7021 7701 7055 7735
rect 7481 7701 7515 7735
rect 7481 7497 7515 7531
rect 4997 7429 5031 7463
rect 2329 7361 2363 7395
rect 4445 7361 4479 7395
rect 4537 7361 4571 7395
rect 5365 7361 5399 7395
rect 7205 7361 7239 7395
rect 2605 7293 2639 7327
rect 4353 7293 4387 7327
rect 5181 7293 5215 7327
rect 5273 7293 5307 7327
rect 6193 7293 6227 7327
rect 6929 7293 6963 7327
rect 4077 7157 4111 7191
rect 4169 7157 4203 7191
rect 5549 7157 5583 7191
rect 6377 7157 6411 7191
rect 4445 6953 4479 6987
rect 5806 6953 5840 6987
rect 7297 6953 7331 6987
rect 5181 6885 5215 6919
rect 3341 6817 3375 6851
rect 4077 6817 4111 6851
rect 5549 6817 5583 6851
rect 3985 6749 4019 6783
rect 4169 6749 4203 6783
rect 4261 6749 4295 6783
rect 4445 6749 4479 6783
rect 4537 6749 4571 6783
rect 4997 6749 5031 6783
rect 5089 6749 5123 6783
rect 5273 6749 5307 6783
rect 7573 6749 7607 6783
rect 3065 6681 3099 6715
rect 3801 6681 3835 6715
rect 5457 6681 5491 6715
rect 1593 6613 1627 6647
rect 4813 6613 4847 6647
rect 7389 6613 7423 6647
rect 2697 6409 2731 6443
rect 3985 6409 4019 6443
rect 5273 6409 5307 6443
rect 6377 6409 6411 6443
rect 7481 6409 7515 6443
rect 1501 6273 1535 6307
rect 1685 6273 1719 6307
rect 2605 6273 2639 6307
rect 2881 6273 2915 6307
rect 3157 6273 3191 6307
rect 4169 6273 4203 6307
rect 5089 6273 5123 6307
rect 6561 6273 6595 6307
rect 6837 6273 6871 6307
rect 7021 6273 7055 6307
rect 7297 6273 7331 6307
rect 2973 6205 3007 6239
rect 3433 6205 3467 6239
rect 3617 6205 3651 6239
rect 3709 6205 3743 6239
rect 3801 6205 3835 6239
rect 4445 6205 4479 6239
rect 4813 6205 4847 6239
rect 6653 6205 6687 6239
rect 6745 6205 6779 6239
rect 3065 6137 3099 6171
rect 2421 6069 2455 6103
rect 4353 6069 4387 6103
rect 4905 6069 4939 6103
rect 2881 5865 2915 5899
rect 3157 5865 3191 5899
rect 5089 5865 5123 5899
rect 3525 5797 3559 5831
rect 2789 5729 2823 5763
rect 2697 5661 2731 5695
rect 3341 5661 3375 5695
rect 3617 5661 3651 5695
rect 7205 5661 7239 5695
rect 3801 5593 3835 5627
rect 3065 5525 3099 5559
rect 7481 5525 7515 5559
rect 4445 5321 4479 5355
rect 3985 5253 4019 5287
rect 1409 5185 1443 5219
rect 3617 5185 3651 5219
rect 3709 5185 3743 5219
rect 4077 5185 4111 5219
rect 4261 5185 4295 5219
rect 5365 5185 5399 5219
rect 5641 5185 5675 5219
rect 3801 5117 3835 5151
rect 5457 5049 5491 5083
rect 1593 4981 1627 5015
rect 4077 4981 4111 5015
rect 5825 4981 5859 5015
rect 2237 4777 2271 4811
rect 4905 4777 4939 4811
rect 2881 4709 2915 4743
rect 2329 4641 2363 4675
rect 3985 4641 4019 4675
rect 4997 4641 5031 4675
rect 2237 4573 2271 4607
rect 2789 4573 2823 4607
rect 2973 4573 3007 4607
rect 3065 4573 3099 4607
rect 4077 4573 4111 4607
rect 4169 4573 4203 4607
rect 4353 4573 4387 4607
rect 4905 4573 4939 4607
rect 5365 4573 5399 4607
rect 7297 4573 7331 4607
rect 3801 4505 3835 4539
rect 5641 4505 5675 4539
rect 2605 4437 2639 4471
rect 3249 4437 3283 4471
rect 4537 4437 4571 4471
rect 5273 4437 5307 4471
rect 7113 4437 7147 4471
rect 7481 4437 7515 4471
rect 4629 4233 4663 4267
rect 6929 4165 6963 4199
rect 1501 4097 1535 4131
rect 1685 4097 1719 4131
rect 1961 4097 1995 4131
rect 3985 4097 4019 4131
rect 4261 4097 4295 4131
rect 4813 4097 4847 4131
rect 4905 4097 4939 4131
rect 5089 4097 5123 4131
rect 5365 4097 5399 4131
rect 5457 4097 5491 4131
rect 5641 4097 5675 4131
rect 6745 4097 6779 4131
rect 7205 4097 7239 4131
rect 2237 4029 2271 4063
rect 3801 4029 3835 4063
rect 6561 4029 6595 4063
rect 6653 4029 6687 4063
rect 7113 4029 7147 4063
rect 7297 4029 7331 4063
rect 3709 3961 3743 3995
rect 4077 3961 4111 3995
rect 4169 3961 4203 3995
rect 4997 3961 5031 3995
rect 5549 3961 5583 3995
rect 6377 3961 6411 3995
rect 1869 3893 1903 3927
rect 5825 3893 5859 3927
rect 4169 3689 4203 3723
rect 4997 3689 5031 3723
rect 5273 3689 5307 3723
rect 1777 3553 1811 3587
rect 4997 3553 5031 3587
rect 5365 3553 5399 3587
rect 5641 3553 5675 3587
rect 4353 3485 4387 3519
rect 4537 3485 4571 3519
rect 4629 3485 4663 3519
rect 4928 3479 4962 3513
rect 7297 3485 7331 3519
rect 2053 3417 2087 3451
rect 3525 3349 3559 3383
rect 7113 3349 7147 3383
rect 7481 3349 7515 3383
rect 5549 3145 5583 3179
rect 6377 3145 6411 3179
rect 4537 3077 4571 3111
rect 1409 3009 1443 3043
rect 5733 3009 5767 3043
rect 6009 3009 6043 3043
rect 6929 3009 6963 3043
rect 7297 3009 7331 3043
rect 1685 2941 1719 2975
rect 5917 2941 5951 2975
rect 3249 2873 3283 2907
rect 7481 2805 7515 2839
rect 3985 2601 4019 2635
rect 4169 2601 4203 2635
rect 3801 2397 3835 2431
rect 3985 2397 4019 2431
rect 7021 2397 7055 2431
rect 7113 2261 7147 2295
<< metal1 >>
rect 1104 8730 7912 8752
rect 1104 8678 2461 8730
rect 2513 8678 2525 8730
rect 2577 8678 2589 8730
rect 2641 8678 2653 8730
rect 2705 8678 2717 8730
rect 2769 8678 4163 8730
rect 4215 8678 4227 8730
rect 4279 8678 4291 8730
rect 4343 8678 4355 8730
rect 4407 8678 4419 8730
rect 4471 8678 5865 8730
rect 5917 8678 5929 8730
rect 5981 8678 5993 8730
rect 6045 8678 6057 8730
rect 6109 8678 6121 8730
rect 6173 8678 7567 8730
rect 7619 8678 7631 8730
rect 7683 8678 7695 8730
rect 7747 8678 7759 8730
rect 7811 8678 7823 8730
rect 7875 8678 7912 8730
rect 1104 8656 7912 8678
rect 6638 8576 6644 8628
rect 6696 8576 6702 8628
rect 1489 8483 1547 8489
rect 1489 8480 1501 8483
rect 204 8452 1501 8480
rect 1489 8449 1501 8452
rect 1535 8449 1547 8483
rect 1489 8443 1547 8449
rect 3605 8483 3663 8489
rect 3605 8449 3617 8483
rect 3651 8480 3663 8483
rect 5074 8480 5080 8492
rect 3651 8452 5080 8480
rect 3651 8449 3663 8452
rect 3605 8443 3663 8449
rect 5074 8440 5080 8452
rect 5132 8440 5138 8492
rect 6733 8483 6791 8489
rect 6733 8449 6745 8483
rect 6779 8480 6791 8483
rect 7374 8480 7380 8492
rect 6779 8452 7380 8480
rect 6779 8449 6791 8452
rect 6733 8443 6791 8449
rect 7374 8440 7380 8452
rect 7432 8440 7438 8492
rect 7466 8372 7472 8424
rect 7524 8372 7530 8424
rect 1673 8347 1731 8353
rect 1673 8313 1685 8347
rect 1719 8344 1731 8347
rect 2866 8344 2872 8356
rect 1719 8316 2872 8344
rect 1719 8313 1731 8316
rect 1673 8307 1731 8313
rect 2866 8304 2872 8316
rect 2924 8304 2930 8356
rect 6917 8347 6975 8353
rect 6917 8313 6929 8347
rect 6963 8344 6975 8347
rect 7282 8344 7288 8356
rect 6963 8316 7288 8344
rect 6963 8313 6975 8316
rect 6917 8307 6975 8313
rect 7282 8304 7288 8316
rect 7340 8304 7346 8356
rect 2314 8236 2320 8288
rect 2372 8236 2378 8288
rect 1104 8186 7912 8208
rect 1104 8134 1801 8186
rect 1853 8134 1865 8186
rect 1917 8134 1929 8186
rect 1981 8134 1993 8186
rect 2045 8134 2057 8186
rect 2109 8134 3503 8186
rect 3555 8134 3567 8186
rect 3619 8134 3631 8186
rect 3683 8134 3695 8186
rect 3747 8134 3759 8186
rect 3811 8134 5205 8186
rect 5257 8134 5269 8186
rect 5321 8134 5333 8186
rect 5385 8134 5397 8186
rect 5449 8134 5461 8186
rect 5513 8134 6907 8186
rect 6959 8134 6971 8186
rect 7023 8134 7035 8186
rect 7087 8134 7099 8186
rect 7151 8134 7163 8186
rect 7215 8134 7912 8186
rect 1104 8112 7912 8134
rect 2314 8032 2320 8084
rect 2372 8072 2378 8084
rect 5169 8075 5227 8081
rect 2372 8044 2774 8072
rect 2372 8032 2378 8044
rect 2746 7936 2774 8044
rect 5169 8041 5181 8075
rect 5215 8072 5227 8075
rect 6822 8072 6828 8084
rect 5215 8044 6828 8072
rect 5215 8041 5227 8044
rect 5169 8035 5227 8041
rect 6822 8032 6828 8044
rect 6880 8032 6886 8084
rect 5261 7939 5319 7945
rect 5261 7936 5273 7939
rect 2746 7908 5273 7936
rect 5261 7905 5273 7908
rect 5307 7936 5319 7939
rect 5534 7936 5540 7948
rect 5307 7908 5540 7936
rect 5307 7905 5319 7908
rect 5261 7899 5319 7905
rect 5534 7896 5540 7908
rect 5592 7896 5598 7948
rect 1489 7871 1547 7877
rect 1489 7868 1501 7871
rect 158 7840 1501 7868
rect 1489 7837 1501 7840
rect 1535 7837 1547 7871
rect 1489 7831 1547 7837
rect 2685 7871 2743 7877
rect 2685 7837 2697 7871
rect 2731 7868 2743 7871
rect 2731 7840 2765 7868
rect 2731 7837 2743 7840
rect 2685 7831 2743 7837
rect 2222 7760 2228 7812
rect 2280 7800 2286 7812
rect 2700 7800 2728 7831
rect 2866 7828 2872 7880
rect 2924 7828 2930 7880
rect 4522 7868 4528 7880
rect 3068 7840 4528 7868
rect 3068 7800 3096 7840
rect 4522 7828 4528 7840
rect 4580 7828 4586 7880
rect 4890 7828 4896 7880
rect 4948 7828 4954 7880
rect 7285 7871 7343 7877
rect 7285 7868 7297 7871
rect 7024 7840 7297 7868
rect 4985 7803 5043 7809
rect 4985 7800 4997 7803
rect 2280 7772 3096 7800
rect 4632 7772 4997 7800
rect 2280 7760 2286 7772
rect 4632 7744 4660 7772
rect 4985 7769 4997 7772
rect 5031 7769 5043 7803
rect 4985 7763 5043 7769
rect 5169 7803 5227 7809
rect 5169 7769 5181 7803
rect 5215 7800 5227 7803
rect 5258 7800 5264 7812
rect 5215 7772 5264 7800
rect 5215 7769 5227 7772
rect 5169 7763 5227 7769
rect 1578 7692 1584 7744
rect 1636 7692 1642 7744
rect 2958 7692 2964 7744
rect 3016 7692 3022 7744
rect 4614 7692 4620 7744
rect 4672 7692 4678 7744
rect 4709 7735 4767 7741
rect 4709 7701 4721 7735
rect 4755 7732 4767 7735
rect 5184 7732 5212 7763
rect 5258 7760 5264 7772
rect 5316 7760 5322 7812
rect 5537 7803 5595 7809
rect 5537 7769 5549 7803
rect 5583 7769 5595 7803
rect 5537 7763 5595 7769
rect 4755 7704 5212 7732
rect 5552 7732 5580 7763
rect 6270 7760 6276 7812
rect 6328 7760 6334 7812
rect 5718 7732 5724 7744
rect 5552 7704 5724 7732
rect 4755 7701 4767 7704
rect 4709 7695 4767 7701
rect 5718 7692 5724 7704
rect 5776 7692 5782 7744
rect 6914 7692 6920 7744
rect 6972 7732 6978 7744
rect 7024 7741 7052 7840
rect 7285 7837 7297 7840
rect 7331 7868 7343 7871
rect 7466 7868 7472 7880
rect 7331 7840 7472 7868
rect 7331 7837 7343 7840
rect 7285 7831 7343 7837
rect 7466 7828 7472 7840
rect 7524 7828 7530 7880
rect 7009 7735 7067 7741
rect 7009 7732 7021 7735
rect 6972 7704 7021 7732
rect 6972 7692 6978 7704
rect 7009 7701 7021 7704
rect 7055 7701 7067 7735
rect 7009 7695 7067 7701
rect 7469 7735 7527 7741
rect 7469 7701 7481 7735
rect 7515 7732 7527 7735
rect 8018 7732 8024 7744
rect 7515 7704 8024 7732
rect 7515 7701 7527 7704
rect 7469 7695 7527 7701
rect 8018 7692 8024 7704
rect 8076 7692 8082 7744
rect 1104 7642 7912 7664
rect 1104 7590 2461 7642
rect 2513 7590 2525 7642
rect 2577 7590 2589 7642
rect 2641 7590 2653 7642
rect 2705 7590 2717 7642
rect 2769 7590 4163 7642
rect 4215 7590 4227 7642
rect 4279 7590 4291 7642
rect 4343 7590 4355 7642
rect 4407 7590 4419 7642
rect 4471 7590 5865 7642
rect 5917 7590 5929 7642
rect 5981 7590 5993 7642
rect 6045 7590 6057 7642
rect 6109 7590 6121 7642
rect 6173 7590 7567 7642
rect 7619 7590 7631 7642
rect 7683 7590 7695 7642
rect 7747 7590 7759 7642
rect 7811 7590 7823 7642
rect 7875 7590 7912 7642
rect 1104 7568 7912 7590
rect 1578 7488 1584 7540
rect 1636 7528 1642 7540
rect 6270 7528 6276 7540
rect 1636 7500 3924 7528
rect 1636 7488 1642 7500
rect 3896 7460 3924 7500
rect 4724 7500 6276 7528
rect 4724 7460 4752 7500
rect 6270 7488 6276 7500
rect 6328 7488 6334 7540
rect 7469 7531 7527 7537
rect 7469 7497 7481 7531
rect 7515 7528 7527 7531
rect 7926 7528 7932 7540
rect 7515 7500 7932 7528
rect 7515 7497 7527 7500
rect 7469 7491 7527 7497
rect 7926 7488 7932 7500
rect 7984 7488 7990 7540
rect 3818 7432 4752 7460
rect 4982 7420 4988 7472
rect 5040 7420 5046 7472
rect 6914 7460 6920 7472
rect 5276 7432 6920 7460
rect 2314 7352 2320 7404
rect 2372 7352 2378 7404
rect 4430 7352 4436 7404
rect 4488 7352 4494 7404
rect 4525 7395 4583 7401
rect 4525 7361 4537 7395
rect 4571 7392 4583 7395
rect 5276 7392 5304 7432
rect 6914 7420 6920 7432
rect 6972 7420 6978 7472
rect 4571 7364 5304 7392
rect 5353 7395 5411 7401
rect 4571 7361 4583 7364
rect 4525 7355 4583 7361
rect 5353 7361 5365 7395
rect 5399 7392 5411 7395
rect 7193 7395 7251 7401
rect 7193 7392 7205 7395
rect 5399 7364 7205 7392
rect 5399 7361 5411 7364
rect 5353 7355 5411 7361
rect 7193 7361 7205 7364
rect 7239 7392 7251 7395
rect 7466 7392 7472 7404
rect 7239 7364 7472 7392
rect 7239 7361 7251 7364
rect 7193 7355 7251 7361
rect 7466 7352 7472 7364
rect 7524 7352 7530 7404
rect 2593 7327 2651 7333
rect 2593 7293 2605 7327
rect 2639 7324 2651 7327
rect 3326 7324 3332 7336
rect 2639 7296 3332 7324
rect 2639 7293 2651 7296
rect 2593 7287 2651 7293
rect 3326 7284 3332 7296
rect 3384 7284 3390 7336
rect 3602 7284 3608 7336
rect 3660 7324 3666 7336
rect 4341 7327 4399 7333
rect 4341 7324 4353 7327
rect 3660 7296 4353 7324
rect 3660 7284 3666 7296
rect 4341 7293 4353 7296
rect 4387 7293 4399 7327
rect 4890 7324 4896 7336
rect 4341 7287 4399 7293
rect 4816 7296 4896 7324
rect 3970 7148 3976 7200
rect 4028 7188 4034 7200
rect 4065 7191 4123 7197
rect 4065 7188 4077 7191
rect 4028 7160 4077 7188
rect 4028 7148 4034 7160
rect 4065 7157 4077 7160
rect 4111 7157 4123 7191
rect 4065 7151 4123 7157
rect 4154 7148 4160 7200
rect 4212 7148 4218 7200
rect 4356 7188 4384 7287
rect 4816 7188 4844 7296
rect 4890 7284 4896 7296
rect 4948 7324 4954 7336
rect 5169 7327 5227 7333
rect 5169 7324 5181 7327
rect 4948 7296 5181 7324
rect 4948 7284 4954 7296
rect 5169 7293 5181 7296
rect 5215 7293 5227 7327
rect 5169 7287 5227 7293
rect 5258 7284 5264 7336
rect 5316 7284 5322 7336
rect 6181 7327 6239 7333
rect 6181 7293 6193 7327
rect 6227 7324 6239 7327
rect 6362 7324 6368 7336
rect 6227 7296 6368 7324
rect 6227 7293 6239 7296
rect 6181 7287 6239 7293
rect 6362 7284 6368 7296
rect 6420 7284 6426 7336
rect 6638 7284 6644 7336
rect 6696 7284 6702 7336
rect 6914 7284 6920 7336
rect 6972 7284 6978 7336
rect 5276 7256 5304 7284
rect 6656 7256 6684 7284
rect 5276 7228 6684 7256
rect 4356 7160 4844 7188
rect 5537 7191 5595 7197
rect 5537 7157 5549 7191
rect 5583 7188 5595 7191
rect 5626 7188 5632 7200
rect 5583 7160 5632 7188
rect 5583 7157 5595 7160
rect 5537 7151 5595 7157
rect 5626 7148 5632 7160
rect 5684 7148 5690 7200
rect 5810 7148 5816 7200
rect 5868 7188 5874 7200
rect 6365 7191 6423 7197
rect 6365 7188 6377 7191
rect 5868 7160 6377 7188
rect 5868 7148 5874 7160
rect 6365 7157 6377 7160
rect 6411 7157 6423 7191
rect 6365 7151 6423 7157
rect 1104 7098 7912 7120
rect 1104 7046 1801 7098
rect 1853 7046 1865 7098
rect 1917 7046 1929 7098
rect 1981 7046 1993 7098
rect 2045 7046 2057 7098
rect 2109 7046 3503 7098
rect 3555 7046 3567 7098
rect 3619 7046 3631 7098
rect 3683 7046 3695 7098
rect 3747 7046 3759 7098
rect 3811 7046 5205 7098
rect 5257 7046 5269 7098
rect 5321 7046 5333 7098
rect 5385 7046 5397 7098
rect 5449 7046 5461 7098
rect 5513 7046 6907 7098
rect 6959 7046 6971 7098
rect 7023 7046 7035 7098
rect 7087 7046 7099 7098
rect 7151 7046 7163 7098
rect 7215 7046 7912 7098
rect 1104 7024 7912 7046
rect 2314 6944 2320 6996
rect 2372 6984 2378 6996
rect 2372 6956 3372 6984
rect 2372 6944 2378 6956
rect 3344 6857 3372 6956
rect 3694 6944 3700 6996
rect 3752 6984 3758 6996
rect 4433 6987 4491 6993
rect 4433 6984 4445 6987
rect 3752 6956 4445 6984
rect 3752 6944 3758 6956
rect 4433 6953 4445 6956
rect 4479 6984 4491 6987
rect 4614 6984 4620 6996
rect 4479 6956 4620 6984
rect 4479 6953 4491 6956
rect 4433 6947 4491 6953
rect 4614 6944 4620 6956
rect 4672 6944 4678 6996
rect 5626 6944 5632 6996
rect 5684 6984 5690 6996
rect 5794 6987 5852 6993
rect 5794 6984 5806 6987
rect 5684 6956 5806 6984
rect 5684 6944 5690 6956
rect 5794 6953 5806 6956
rect 5840 6953 5852 6987
rect 5794 6947 5852 6953
rect 7285 6987 7343 6993
rect 7285 6953 7297 6987
rect 7331 6984 7343 6987
rect 7466 6984 7472 6996
rect 7331 6956 7472 6984
rect 7331 6953 7343 6956
rect 7285 6947 7343 6953
rect 7466 6944 7472 6956
rect 7524 6944 7530 6996
rect 4154 6876 4160 6928
rect 4212 6876 4218 6928
rect 4982 6876 4988 6928
rect 5040 6916 5046 6928
rect 5169 6919 5227 6925
rect 5169 6916 5181 6919
rect 5040 6888 5181 6916
rect 5040 6876 5046 6888
rect 5169 6885 5181 6888
rect 5215 6885 5227 6919
rect 5169 6879 5227 6885
rect 5460 6888 5672 6916
rect 3329 6851 3387 6857
rect 3329 6817 3341 6851
rect 3375 6817 3387 6851
rect 3329 6811 3387 6817
rect 4065 6851 4123 6857
rect 4065 6817 4077 6851
rect 4111 6848 4123 6851
rect 4172 6848 4200 6876
rect 5460 6848 5488 6888
rect 4111 6820 4200 6848
rect 4448 6820 5488 6848
rect 4111 6817 4123 6820
rect 4065 6811 4123 6817
rect 1578 6740 1584 6792
rect 1636 6780 1642 6792
rect 1636 6752 1978 6780
rect 1636 6740 1642 6752
rect 3878 6740 3884 6792
rect 3936 6780 3942 6792
rect 4448 6789 4476 6820
rect 5534 6808 5540 6860
rect 5592 6808 5598 6860
rect 5644 6848 5672 6888
rect 5810 6848 5816 6860
rect 5644 6820 5816 6848
rect 5810 6808 5816 6820
rect 5868 6808 5874 6860
rect 3973 6783 4031 6789
rect 3973 6780 3985 6783
rect 3936 6752 3985 6780
rect 3936 6740 3942 6752
rect 3973 6749 3985 6752
rect 4019 6749 4031 6783
rect 3973 6743 4031 6749
rect 4157 6783 4215 6789
rect 4157 6749 4169 6783
rect 4203 6749 4215 6783
rect 4157 6743 4215 6749
rect 4249 6783 4307 6789
rect 4249 6749 4261 6783
rect 4295 6749 4307 6783
rect 4249 6743 4307 6749
rect 4433 6783 4491 6789
rect 4433 6749 4445 6783
rect 4479 6749 4491 6783
rect 4433 6743 4491 6749
rect 3050 6672 3056 6724
rect 3108 6672 3114 6724
rect 3326 6672 3332 6724
rect 3384 6712 3390 6724
rect 3789 6715 3847 6721
rect 3789 6712 3801 6715
rect 3384 6684 3801 6712
rect 3384 6672 3390 6684
rect 3789 6681 3801 6684
rect 3835 6681 3847 6715
rect 3789 6675 3847 6681
rect 4062 6672 4068 6724
rect 4120 6712 4126 6724
rect 4172 6712 4200 6743
rect 4120 6684 4200 6712
rect 4120 6672 4126 6684
rect 1578 6604 1584 6656
rect 1636 6604 1642 6656
rect 2866 6604 2872 6656
rect 2924 6644 2930 6656
rect 3694 6644 3700 6656
rect 2924 6616 3700 6644
rect 2924 6604 2930 6616
rect 3694 6604 3700 6616
rect 3752 6604 3758 6656
rect 4264 6644 4292 6743
rect 4522 6740 4528 6792
rect 4580 6740 4586 6792
rect 4985 6783 5043 6789
rect 4985 6780 4997 6783
rect 4816 6752 4997 6780
rect 4522 6644 4528 6656
rect 4264 6616 4528 6644
rect 4522 6604 4528 6616
rect 4580 6604 4586 6656
rect 4816 6653 4844 6752
rect 4985 6749 4997 6752
rect 5031 6749 5043 6783
rect 4985 6743 5043 6749
rect 5077 6783 5135 6789
rect 5077 6749 5089 6783
rect 5123 6780 5135 6783
rect 5166 6780 5172 6792
rect 5123 6752 5172 6780
rect 5123 6749 5135 6752
rect 5077 6743 5135 6749
rect 5166 6740 5172 6752
rect 5224 6740 5230 6792
rect 5261 6783 5319 6789
rect 5261 6749 5273 6783
rect 5307 6749 5319 6783
rect 7484 6780 7512 6944
rect 7561 6783 7619 6789
rect 7561 6780 7573 6783
rect 7484 6752 7573 6780
rect 5261 6743 5319 6749
rect 7561 6749 7573 6752
rect 7607 6749 7619 6783
rect 7561 6743 7619 6749
rect 5276 6712 5304 6743
rect 4908 6684 5304 6712
rect 5445 6715 5503 6721
rect 4908 6656 4936 6684
rect 5445 6681 5457 6715
rect 5491 6712 5503 6715
rect 5718 6712 5724 6724
rect 5491 6684 5724 6712
rect 5491 6681 5503 6684
rect 5445 6675 5503 6681
rect 5718 6672 5724 6684
rect 5776 6672 5782 6724
rect 6270 6672 6276 6724
rect 6328 6672 6334 6724
rect 4801 6647 4859 6653
rect 4801 6613 4813 6647
rect 4847 6613 4859 6647
rect 4801 6607 4859 6613
rect 4890 6604 4896 6656
rect 4948 6604 4954 6656
rect 7374 6604 7380 6656
rect 7432 6604 7438 6656
rect 1104 6554 7912 6576
rect 1104 6502 2461 6554
rect 2513 6502 2525 6554
rect 2577 6502 2589 6554
rect 2641 6502 2653 6554
rect 2705 6502 2717 6554
rect 2769 6502 4163 6554
rect 4215 6502 4227 6554
rect 4279 6502 4291 6554
rect 4343 6502 4355 6554
rect 4407 6502 4419 6554
rect 4471 6502 5865 6554
rect 5917 6502 5929 6554
rect 5981 6502 5993 6554
rect 6045 6502 6057 6554
rect 6109 6502 6121 6554
rect 6173 6502 7567 6554
rect 7619 6502 7631 6554
rect 7683 6502 7695 6554
rect 7747 6502 7759 6554
rect 7811 6502 7823 6554
rect 7875 6502 7912 6554
rect 1104 6480 7912 6502
rect 2685 6443 2743 6449
rect 2685 6409 2697 6443
rect 2731 6440 2743 6443
rect 3050 6440 3056 6452
rect 2731 6412 3056 6440
rect 2731 6409 2743 6412
rect 2685 6403 2743 6409
rect 3050 6400 3056 6412
rect 3108 6400 3114 6452
rect 3973 6443 4031 6449
rect 3973 6409 3985 6443
rect 4019 6440 4031 6443
rect 4062 6440 4068 6452
rect 4019 6412 4068 6440
rect 4019 6409 4031 6412
rect 3973 6403 4031 6409
rect 4062 6400 4068 6412
rect 4120 6400 4126 6452
rect 5166 6400 5172 6452
rect 5224 6440 5230 6452
rect 5261 6443 5319 6449
rect 5261 6440 5273 6443
rect 5224 6412 5273 6440
rect 5224 6400 5230 6412
rect 5261 6409 5273 6412
rect 5307 6409 5319 6443
rect 5261 6403 5319 6409
rect 6362 6400 6368 6452
rect 6420 6400 6426 6452
rect 7469 6443 7527 6449
rect 6472 6412 7328 6440
rect 2958 6372 2964 6384
rect 2884 6344 2964 6372
rect 1489 6307 1547 6313
rect 1489 6304 1501 6307
rect 472 6276 1501 6304
rect 1489 6273 1501 6276
rect 1535 6273 1547 6307
rect 1489 6267 1547 6273
rect 1673 6307 1731 6313
rect 1673 6273 1685 6307
rect 1719 6304 1731 6307
rect 2222 6304 2228 6316
rect 1719 6276 2228 6304
rect 1719 6273 1731 6276
rect 1673 6267 1731 6273
rect 2222 6264 2228 6276
rect 2280 6304 2286 6316
rect 2590 6304 2596 6316
rect 2280 6276 2596 6304
rect 2280 6264 2286 6276
rect 2590 6264 2596 6276
rect 2648 6264 2654 6316
rect 2884 6313 2912 6344
rect 2958 6332 2964 6344
rect 3016 6372 3022 6384
rect 3878 6372 3884 6384
rect 3016 6344 3884 6372
rect 3016 6332 3022 6344
rect 3878 6332 3884 6344
rect 3936 6372 3942 6384
rect 4890 6372 4896 6384
rect 3936 6344 4896 6372
rect 3936 6332 3942 6344
rect 4890 6332 4896 6344
rect 4948 6332 4954 6384
rect 2869 6307 2927 6313
rect 2869 6273 2881 6307
rect 2915 6273 2927 6307
rect 2869 6267 2927 6273
rect 3142 6264 3148 6316
rect 3200 6264 3206 6316
rect 4157 6307 4215 6313
rect 4157 6273 4169 6307
rect 4203 6304 4215 6307
rect 4246 6304 4252 6316
rect 4203 6276 4252 6304
rect 4203 6273 4215 6276
rect 4157 6267 4215 6273
rect 4246 6264 4252 6276
rect 4304 6264 4310 6316
rect 5077 6307 5135 6313
rect 5077 6304 5089 6307
rect 4356 6276 5089 6304
rect 2961 6239 3019 6245
rect 2961 6205 2973 6239
rect 3007 6236 3019 6239
rect 3421 6239 3479 6245
rect 3421 6236 3433 6239
rect 3007 6208 3433 6236
rect 3007 6205 3019 6208
rect 2961 6199 3019 6205
rect 3421 6205 3433 6208
rect 3467 6205 3479 6239
rect 3421 6199 3479 6205
rect 3510 6196 3516 6248
rect 3568 6236 3574 6248
rect 3605 6239 3663 6245
rect 3605 6236 3617 6239
rect 3568 6208 3617 6236
rect 3568 6196 3574 6208
rect 3605 6205 3617 6208
rect 3651 6205 3663 6239
rect 3605 6199 3663 6205
rect 3697 6239 3755 6245
rect 3697 6205 3709 6239
rect 3743 6205 3755 6239
rect 3697 6199 3755 6205
rect 3789 6239 3847 6245
rect 3789 6205 3801 6239
rect 3835 6236 3847 6239
rect 3970 6236 3976 6248
rect 3835 6208 3976 6236
rect 3835 6205 3847 6208
rect 3789 6199 3847 6205
rect 3050 6128 3056 6180
rect 3108 6128 3114 6180
rect 3712 6168 3740 6199
rect 3970 6196 3976 6208
rect 4028 6236 4034 6248
rect 4356 6236 4384 6276
rect 5077 6273 5089 6276
rect 5123 6304 5135 6307
rect 6472 6304 6500 6412
rect 6638 6332 6644 6384
rect 6696 6332 6702 6384
rect 7098 6372 7104 6384
rect 6840 6344 7104 6372
rect 5123 6276 6500 6304
rect 6549 6307 6607 6313
rect 5123 6273 5135 6276
rect 5077 6267 5135 6273
rect 6549 6273 6561 6307
rect 6595 6304 6607 6307
rect 6656 6304 6684 6332
rect 6840 6313 6868 6344
rect 7098 6332 7104 6344
rect 7156 6332 7162 6384
rect 6595 6276 6684 6304
rect 6825 6307 6883 6313
rect 6595 6273 6607 6276
rect 6549 6267 6607 6273
rect 6825 6273 6837 6307
rect 6871 6273 6883 6307
rect 6825 6267 6883 6273
rect 6914 6264 6920 6316
rect 6972 6304 6978 6316
rect 7300 6313 7328 6412
rect 7469 6409 7481 6443
rect 7515 6440 7527 6443
rect 8018 6440 8024 6452
rect 7515 6412 8024 6440
rect 7515 6409 7527 6412
rect 7469 6403 7527 6409
rect 8018 6400 8024 6412
rect 8076 6400 8082 6452
rect 7009 6307 7067 6313
rect 7009 6304 7021 6307
rect 6972 6276 7021 6304
rect 6972 6264 6978 6276
rect 7009 6273 7021 6276
rect 7055 6273 7067 6307
rect 7009 6267 7067 6273
rect 7285 6307 7343 6313
rect 7285 6273 7297 6307
rect 7331 6273 7343 6307
rect 7285 6267 7343 6273
rect 7466 6264 7472 6316
rect 7524 6264 7530 6316
rect 4028 6208 4384 6236
rect 4433 6239 4491 6245
rect 4028 6196 4034 6208
rect 4433 6205 4445 6239
rect 4479 6236 4491 6239
rect 4798 6236 4804 6248
rect 4479 6208 4804 6236
rect 4479 6205 4491 6208
rect 4433 6199 4491 6205
rect 3878 6168 3884 6180
rect 3712 6140 3884 6168
rect 3878 6128 3884 6140
rect 3936 6128 3942 6180
rect 4448 6168 4476 6199
rect 4798 6196 4804 6208
rect 4856 6196 4862 6248
rect 4890 6196 4896 6248
rect 4948 6236 4954 6248
rect 6641 6239 6699 6245
rect 6641 6236 6653 6239
rect 4948 6208 6653 6236
rect 4948 6196 4954 6208
rect 6641 6205 6653 6208
rect 6687 6205 6699 6239
rect 6641 6199 6699 6205
rect 6733 6239 6791 6245
rect 6733 6205 6745 6239
rect 6779 6236 6791 6239
rect 7484 6236 7512 6264
rect 6779 6208 7512 6236
rect 6779 6205 6791 6208
rect 6733 6199 6791 6205
rect 4264 6140 4476 6168
rect 2314 6060 2320 6112
rect 2372 6100 2378 6112
rect 2409 6103 2467 6109
rect 2409 6100 2421 6103
rect 2372 6072 2421 6100
rect 2372 6060 2378 6072
rect 2409 6069 2421 6072
rect 2455 6100 2467 6103
rect 4264 6100 4292 6140
rect 2455 6072 4292 6100
rect 2455 6069 2467 6072
rect 2409 6063 2467 6069
rect 4338 6060 4344 6112
rect 4396 6100 4402 6112
rect 4893 6103 4951 6109
rect 4893 6100 4905 6103
rect 4396 6072 4905 6100
rect 4396 6060 4402 6072
rect 4893 6069 4905 6072
rect 4939 6069 4951 6103
rect 4893 6063 4951 6069
rect 1104 6010 7912 6032
rect 1104 5958 1801 6010
rect 1853 5958 1865 6010
rect 1917 5958 1929 6010
rect 1981 5958 1993 6010
rect 2045 5958 2057 6010
rect 2109 5958 3503 6010
rect 3555 5958 3567 6010
rect 3619 5958 3631 6010
rect 3683 5958 3695 6010
rect 3747 5958 3759 6010
rect 3811 5958 5205 6010
rect 5257 5958 5269 6010
rect 5321 5958 5333 6010
rect 5385 5958 5397 6010
rect 5449 5958 5461 6010
rect 5513 5958 6907 6010
rect 6959 5958 6971 6010
rect 7023 5958 7035 6010
rect 7087 5958 7099 6010
rect 7151 5958 7163 6010
rect 7215 5958 7912 6010
rect 1104 5936 7912 5958
rect 2222 5856 2228 5908
rect 2280 5896 2286 5908
rect 2866 5896 2872 5908
rect 2280 5868 2872 5896
rect 2280 5856 2286 5868
rect 2866 5856 2872 5868
rect 2924 5856 2930 5908
rect 3050 5856 3056 5908
rect 3108 5896 3114 5908
rect 3145 5899 3203 5905
rect 3145 5896 3157 5899
rect 3108 5868 3157 5896
rect 3108 5856 3114 5868
rect 3145 5865 3157 5868
rect 3191 5865 3203 5899
rect 3145 5859 3203 5865
rect 5074 5856 5080 5908
rect 5132 5856 5138 5908
rect 3513 5831 3571 5837
rect 3513 5797 3525 5831
rect 3559 5828 3571 5831
rect 4338 5828 4344 5840
rect 3559 5800 4344 5828
rect 3559 5797 3571 5800
rect 3513 5791 3571 5797
rect 4338 5788 4344 5800
rect 4396 5828 4402 5840
rect 4396 5800 4752 5828
rect 4396 5788 4402 5800
rect 4724 5772 4752 5800
rect 2590 5720 2596 5772
rect 2648 5760 2654 5772
rect 2777 5763 2835 5769
rect 2777 5760 2789 5763
rect 2648 5732 2789 5760
rect 2648 5720 2654 5732
rect 2777 5729 2789 5732
rect 2823 5729 2835 5763
rect 2777 5723 2835 5729
rect 4706 5720 4712 5772
rect 4764 5720 4770 5772
rect 1578 5652 1584 5704
rect 1636 5692 1642 5704
rect 2685 5695 2743 5701
rect 2685 5692 2697 5695
rect 1636 5664 2697 5692
rect 1636 5652 1642 5664
rect 2685 5661 2697 5664
rect 2731 5661 2743 5695
rect 2685 5655 2743 5661
rect 2700 5556 2728 5655
rect 3326 5652 3332 5704
rect 3384 5652 3390 5704
rect 3510 5652 3516 5704
rect 3568 5692 3574 5704
rect 3605 5695 3663 5701
rect 3605 5692 3617 5695
rect 3568 5664 3617 5692
rect 3568 5652 3574 5664
rect 3605 5661 3617 5664
rect 3651 5661 3663 5695
rect 3605 5655 3663 5661
rect 3694 5652 3700 5704
rect 3752 5692 3758 5704
rect 4246 5692 4252 5704
rect 3752 5664 4252 5692
rect 3752 5652 3758 5664
rect 4246 5652 4252 5664
rect 4304 5692 4310 5704
rect 7193 5695 7251 5701
rect 7193 5692 7205 5695
rect 4304 5664 7205 5692
rect 4304 5652 4310 5664
rect 7193 5661 7205 5664
rect 7239 5661 7251 5695
rect 7193 5655 7251 5661
rect 2866 5584 2872 5636
rect 2924 5624 2930 5636
rect 3789 5627 3847 5633
rect 3789 5624 3801 5627
rect 2924 5596 3801 5624
rect 2924 5584 2930 5596
rect 3789 5593 3801 5596
rect 3835 5593 3847 5627
rect 3789 5587 3847 5593
rect 2958 5556 2964 5568
rect 2700 5528 2964 5556
rect 2958 5516 2964 5528
rect 3016 5516 3022 5568
rect 3053 5559 3111 5565
rect 3053 5525 3065 5559
rect 3099 5556 3111 5559
rect 3142 5556 3148 5568
rect 3099 5528 3148 5556
rect 3099 5525 3111 5528
rect 3053 5519 3111 5525
rect 3142 5516 3148 5528
rect 3200 5516 3206 5568
rect 7469 5559 7527 5565
rect 7469 5525 7481 5559
rect 7515 5556 7527 5559
rect 8018 5556 8024 5568
rect 7515 5528 8024 5556
rect 7515 5525 7527 5528
rect 7469 5519 7527 5525
rect 8018 5516 8024 5528
rect 8076 5516 8082 5568
rect 1104 5466 7912 5488
rect 1104 5414 2461 5466
rect 2513 5414 2525 5466
rect 2577 5414 2589 5466
rect 2641 5414 2653 5466
rect 2705 5414 2717 5466
rect 2769 5414 4163 5466
rect 4215 5414 4227 5466
rect 4279 5414 4291 5466
rect 4343 5414 4355 5466
rect 4407 5414 4419 5466
rect 4471 5414 5865 5466
rect 5917 5414 5929 5466
rect 5981 5414 5993 5466
rect 6045 5414 6057 5466
rect 6109 5414 6121 5466
rect 6173 5414 7567 5466
rect 7619 5414 7631 5466
rect 7683 5414 7695 5466
rect 7747 5414 7759 5466
rect 7811 5414 7823 5466
rect 7875 5414 7912 5466
rect 1104 5392 7912 5414
rect 2314 5312 2320 5364
rect 2372 5352 2378 5364
rect 3510 5352 3516 5364
rect 2372 5324 3516 5352
rect 2372 5312 2378 5324
rect 3510 5312 3516 5324
rect 3568 5312 3574 5364
rect 3694 5312 3700 5364
rect 3752 5312 3758 5364
rect 4433 5355 4491 5361
rect 4433 5321 4445 5355
rect 4479 5352 4491 5355
rect 4522 5352 4528 5364
rect 4479 5324 4528 5352
rect 4479 5321 4491 5324
rect 4433 5315 4491 5321
rect 4522 5312 4528 5324
rect 4580 5312 4586 5364
rect 2958 5244 2964 5296
rect 3016 5284 3022 5296
rect 3712 5284 3740 5312
rect 3016 5256 3740 5284
rect 3973 5287 4031 5293
rect 3016 5244 3022 5256
rect 3620 5225 3648 5256
rect 3973 5253 3985 5287
rect 4019 5284 4031 5287
rect 4154 5284 4160 5296
rect 4019 5256 4160 5284
rect 4019 5253 4031 5256
rect 3973 5247 4031 5253
rect 4154 5244 4160 5256
rect 4212 5244 4218 5296
rect 1397 5219 1455 5225
rect 1397 5216 1409 5219
rect 518 5188 1409 5216
rect 1397 5185 1409 5188
rect 1443 5185 1455 5219
rect 1397 5179 1455 5185
rect 3605 5219 3663 5225
rect 3605 5185 3617 5219
rect 3651 5185 3663 5219
rect 3605 5179 3663 5185
rect 3697 5219 3755 5225
rect 3697 5185 3709 5219
rect 3743 5216 3755 5219
rect 3878 5216 3884 5228
rect 3743 5188 3884 5216
rect 3743 5185 3755 5188
rect 3697 5179 3755 5185
rect 3878 5176 3884 5188
rect 3936 5176 3942 5228
rect 4062 5176 4068 5228
rect 4120 5176 4126 5228
rect 4249 5219 4307 5225
rect 4249 5185 4261 5219
rect 4295 5216 4307 5219
rect 4614 5216 4620 5228
rect 4295 5188 4620 5216
rect 4295 5185 4307 5188
rect 4249 5179 4307 5185
rect 4614 5176 4620 5188
rect 4672 5176 4678 5228
rect 4798 5176 4804 5228
rect 4856 5216 4862 5228
rect 5353 5219 5411 5225
rect 5353 5216 5365 5219
rect 4856 5188 5365 5216
rect 4856 5176 4862 5188
rect 5353 5185 5365 5188
rect 5399 5185 5411 5219
rect 5353 5179 5411 5185
rect 5629 5219 5687 5225
rect 5629 5185 5641 5219
rect 5675 5216 5687 5219
rect 7374 5216 7380 5228
rect 5675 5188 7380 5216
rect 5675 5185 5687 5188
rect 5629 5179 5687 5185
rect 7374 5176 7380 5188
rect 7432 5176 7438 5228
rect 3418 5108 3424 5160
rect 3476 5148 3482 5160
rect 3789 5151 3847 5157
rect 3789 5148 3801 5151
rect 3476 5120 3801 5148
rect 3476 5108 3482 5120
rect 3789 5117 3801 5120
rect 3835 5117 3847 5151
rect 3789 5111 3847 5117
rect 3804 5080 3832 5111
rect 3970 5108 3976 5160
rect 4028 5148 4034 5160
rect 6270 5148 6276 5160
rect 4028 5120 6276 5148
rect 4028 5108 4034 5120
rect 6270 5108 6276 5120
rect 6328 5108 6334 5160
rect 4430 5080 4436 5092
rect 3804 5052 4436 5080
rect 4430 5040 4436 5052
rect 4488 5080 4494 5092
rect 5445 5083 5503 5089
rect 5445 5080 5457 5083
rect 4488 5052 5457 5080
rect 4488 5040 4494 5052
rect 5445 5049 5457 5052
rect 5491 5080 5503 5083
rect 5491 5052 6592 5080
rect 5491 5049 5503 5052
rect 5445 5043 5503 5049
rect 6564 5024 6592 5052
rect 1578 4972 1584 5024
rect 1636 4972 1642 5024
rect 2222 4972 2228 5024
rect 2280 5012 2286 5024
rect 4065 5015 4123 5021
rect 4065 5012 4077 5015
rect 2280 4984 4077 5012
rect 2280 4972 2286 4984
rect 4065 4981 4077 4984
rect 4111 5012 4123 5015
rect 4890 5012 4896 5024
rect 4111 4984 4896 5012
rect 4111 4981 4123 4984
rect 4065 4975 4123 4981
rect 4890 4972 4896 4984
rect 4948 4972 4954 5024
rect 5534 4972 5540 5024
rect 5592 5012 5598 5024
rect 5813 5015 5871 5021
rect 5813 5012 5825 5015
rect 5592 4984 5825 5012
rect 5592 4972 5598 4984
rect 5813 4981 5825 4984
rect 5859 4981 5871 5015
rect 5813 4975 5871 4981
rect 6546 4972 6552 5024
rect 6604 4972 6610 5024
rect 1104 4922 7912 4944
rect 1104 4870 1801 4922
rect 1853 4870 1865 4922
rect 1917 4870 1929 4922
rect 1981 4870 1993 4922
rect 2045 4870 2057 4922
rect 2109 4870 3503 4922
rect 3555 4870 3567 4922
rect 3619 4870 3631 4922
rect 3683 4870 3695 4922
rect 3747 4870 3759 4922
rect 3811 4870 5205 4922
rect 5257 4870 5269 4922
rect 5321 4870 5333 4922
rect 5385 4870 5397 4922
rect 5449 4870 5461 4922
rect 5513 4870 6907 4922
rect 6959 4870 6971 4922
rect 7023 4870 7035 4922
rect 7087 4870 7099 4922
rect 7151 4870 7163 4922
rect 7215 4870 7912 4922
rect 1104 4848 7912 4870
rect 2222 4768 2228 4820
rect 2280 4768 2286 4820
rect 4890 4768 4896 4820
rect 4948 4768 4954 4820
rect 2869 4743 2927 4749
rect 2240 4712 2774 4740
rect 2240 4613 2268 4712
rect 2314 4632 2320 4684
rect 2372 4632 2378 4684
rect 2746 4672 2774 4712
rect 2869 4709 2881 4743
rect 2915 4740 2927 4743
rect 2958 4740 2964 4752
rect 2915 4712 2964 4740
rect 2915 4709 2927 4712
rect 2869 4703 2927 4709
rect 2958 4700 2964 4712
rect 3016 4700 3022 4752
rect 3418 4700 3424 4752
rect 3476 4700 3482 4752
rect 4430 4740 4436 4752
rect 3988 4712 4436 4740
rect 3436 4672 3464 4700
rect 3988 4681 4016 4712
rect 4430 4700 4436 4712
rect 4488 4700 4494 4752
rect 4724 4712 5120 4740
rect 2746 4644 3464 4672
rect 3973 4675 4031 4681
rect 3973 4641 3985 4675
rect 4019 4641 4031 4675
rect 4724 4672 4752 4712
rect 3973 4635 4031 4641
rect 4080 4644 4752 4672
rect 2225 4607 2283 4613
rect 2225 4573 2237 4607
rect 2271 4573 2283 4607
rect 2777 4607 2835 4613
rect 2777 4604 2789 4607
rect 2225 4567 2283 4573
rect 2608 4576 2789 4604
rect 2608 4477 2636 4576
rect 2777 4573 2789 4576
rect 2823 4573 2835 4607
rect 2777 4567 2835 4573
rect 2961 4607 3019 4613
rect 2961 4573 2973 4607
rect 3007 4573 3019 4607
rect 2961 4567 3019 4573
rect 3053 4607 3111 4613
rect 3053 4573 3065 4607
rect 3099 4604 3111 4607
rect 3099 4576 3832 4604
rect 3099 4573 3111 4576
rect 3053 4567 3111 4573
rect 2976 4536 3004 4567
rect 3142 4536 3148 4548
rect 2976 4508 3148 4536
rect 3142 4496 3148 4508
rect 3200 4496 3206 4548
rect 3804 4545 3832 4576
rect 3878 4564 3884 4616
rect 3936 4604 3942 4616
rect 4080 4613 4108 4644
rect 4798 4632 4804 4684
rect 4856 4672 4862 4684
rect 4985 4675 5043 4681
rect 4985 4672 4997 4675
rect 4856 4644 4997 4672
rect 4856 4632 4862 4644
rect 4985 4641 4997 4644
rect 5031 4641 5043 4675
rect 5092 4672 5120 4712
rect 6638 4672 6644 4684
rect 5092 4644 6644 4672
rect 4985 4635 5043 4641
rect 6638 4632 6644 4644
rect 6696 4632 6702 4684
rect 6822 4632 6828 4684
rect 6880 4672 6886 4684
rect 6880 4644 7328 4672
rect 6880 4632 6886 4644
rect 4065 4607 4123 4613
rect 4065 4604 4077 4607
rect 3936 4576 4077 4604
rect 3936 4564 3942 4576
rect 4065 4573 4077 4576
rect 4111 4573 4123 4607
rect 4065 4567 4123 4573
rect 4157 4607 4215 4613
rect 4157 4573 4169 4607
rect 4203 4573 4215 4607
rect 4157 4567 4215 4573
rect 4341 4607 4399 4613
rect 4341 4573 4353 4607
rect 4387 4604 4399 4607
rect 4522 4604 4528 4616
rect 4387 4576 4528 4604
rect 4387 4573 4399 4576
rect 4341 4567 4399 4573
rect 3789 4539 3847 4545
rect 3789 4505 3801 4539
rect 3835 4505 3847 4539
rect 4172 4536 4200 4567
rect 4522 4564 4528 4576
rect 4580 4564 4586 4616
rect 4893 4607 4951 4613
rect 4893 4573 4905 4607
rect 4939 4573 4951 4607
rect 4893 4567 4951 4573
rect 4908 4536 4936 4567
rect 5074 4564 5080 4616
rect 5132 4604 5138 4616
rect 7300 4613 7328 4644
rect 5353 4607 5411 4613
rect 5353 4604 5365 4607
rect 5132 4576 5365 4604
rect 5132 4564 5138 4576
rect 5353 4573 5365 4576
rect 5399 4573 5411 4607
rect 5353 4567 5411 4573
rect 7285 4607 7343 4613
rect 7285 4573 7297 4607
rect 7331 4573 7343 4607
rect 7285 4567 7343 4573
rect 4172 4508 5396 4536
rect 3789 4499 3847 4505
rect 2593 4471 2651 4477
rect 2593 4437 2605 4471
rect 2639 4437 2651 4471
rect 2593 4431 2651 4437
rect 3050 4428 3056 4480
rect 3108 4468 3114 4480
rect 3237 4471 3295 4477
rect 3237 4468 3249 4471
rect 3108 4440 3249 4468
rect 3108 4428 3114 4440
rect 3237 4437 3249 4440
rect 3283 4437 3295 4471
rect 3237 4431 3295 4437
rect 3970 4428 3976 4480
rect 4028 4468 4034 4480
rect 4154 4468 4160 4480
rect 4028 4440 4160 4468
rect 4028 4428 4034 4440
rect 4154 4428 4160 4440
rect 4212 4428 4218 4480
rect 4430 4428 4436 4480
rect 4488 4468 4494 4480
rect 4525 4471 4583 4477
rect 4525 4468 4537 4471
rect 4488 4440 4537 4468
rect 4488 4428 4494 4440
rect 4525 4437 4537 4440
rect 4571 4437 4583 4471
rect 4525 4431 4583 4437
rect 4706 4428 4712 4480
rect 4764 4468 4770 4480
rect 4890 4468 4896 4480
rect 4764 4440 4896 4468
rect 4764 4428 4770 4440
rect 4890 4428 4896 4440
rect 4948 4428 4954 4480
rect 5258 4428 5264 4480
rect 5316 4428 5322 4480
rect 5368 4468 5396 4508
rect 5626 4496 5632 4548
rect 5684 4496 5690 4548
rect 6270 4496 6276 4548
rect 6328 4496 6334 4548
rect 7101 4471 7159 4477
rect 7101 4468 7113 4471
rect 5368 4440 7113 4468
rect 7101 4437 7113 4440
rect 7147 4468 7159 4471
rect 7374 4468 7380 4480
rect 7147 4440 7380 4468
rect 7147 4437 7159 4440
rect 7101 4431 7159 4437
rect 7374 4428 7380 4440
rect 7432 4428 7438 4480
rect 7469 4471 7527 4477
rect 7469 4437 7481 4471
rect 7515 4468 7527 4471
rect 8018 4468 8024 4480
rect 7515 4440 8024 4468
rect 7515 4437 7527 4440
rect 7469 4431 7527 4437
rect 8018 4428 8024 4440
rect 8076 4428 8082 4480
rect 1104 4378 7912 4400
rect 1104 4326 2461 4378
rect 2513 4326 2525 4378
rect 2577 4326 2589 4378
rect 2641 4326 2653 4378
rect 2705 4326 2717 4378
rect 2769 4326 4163 4378
rect 4215 4326 4227 4378
rect 4279 4326 4291 4378
rect 4343 4326 4355 4378
rect 4407 4326 4419 4378
rect 4471 4326 5865 4378
rect 5917 4326 5929 4378
rect 5981 4326 5993 4378
rect 6045 4326 6057 4378
rect 6109 4326 6121 4378
rect 6173 4326 7567 4378
rect 7619 4326 7631 4378
rect 7683 4326 7695 4378
rect 7747 4326 7759 4378
rect 7811 4326 7823 4378
rect 7875 4326 7912 4378
rect 1104 4304 7912 4326
rect 1578 4224 1584 4276
rect 1636 4224 1642 4276
rect 2222 4264 2228 4276
rect 1872 4236 2228 4264
rect 1489 4131 1547 4137
rect 1489 4097 1501 4131
rect 1535 4097 1547 4131
rect 1596 4128 1624 4224
rect 1673 4131 1731 4137
rect 1673 4128 1685 4131
rect 1596 4100 1685 4128
rect 1489 4091 1547 4097
rect 1673 4097 1685 4100
rect 1719 4097 1731 4131
rect 1673 4091 1731 4097
rect 1504 4060 1532 4091
rect 1872 4060 1900 4236
rect 2222 4224 2228 4236
rect 2280 4224 2286 4276
rect 3142 4224 3148 4276
rect 3200 4264 3206 4276
rect 4617 4267 4675 4273
rect 3200 4236 4016 4264
rect 3200 4224 3206 4236
rect 2314 4196 2320 4208
rect 1964 4168 2320 4196
rect 1964 4137 1992 4168
rect 2314 4156 2320 4168
rect 2372 4156 2378 4208
rect 3988 4196 4016 4236
rect 4617 4233 4629 4267
rect 4663 4264 4675 4267
rect 5626 4264 5632 4276
rect 4663 4236 5632 4264
rect 4663 4233 4675 4236
rect 4617 4227 4675 4233
rect 5626 4224 5632 4236
rect 5684 4224 5690 4276
rect 4430 4196 4436 4208
rect 3988 4168 4436 4196
rect 1949 4131 2007 4137
rect 1949 4097 1961 4131
rect 1995 4097 2007 4131
rect 3878 4128 3884 4140
rect 3358 4100 3884 4128
rect 1949 4091 2007 4097
rect 3878 4088 3884 4100
rect 3936 4088 3942 4140
rect 3988 4137 4016 4168
rect 4430 4156 4436 4168
rect 4488 4196 4494 4208
rect 6917 4199 6975 4205
rect 6917 4196 6929 4199
rect 4488 4168 4844 4196
rect 4488 4156 4494 4168
rect 3973 4131 4031 4137
rect 3973 4097 3985 4131
rect 4019 4097 4031 4131
rect 3973 4091 4031 4097
rect 4249 4131 4307 4137
rect 4249 4097 4261 4131
rect 4295 4128 4307 4131
rect 4614 4128 4620 4140
rect 4295 4100 4620 4128
rect 4295 4097 4307 4100
rect 4249 4091 4307 4097
rect 4614 4088 4620 4100
rect 4672 4088 4678 4140
rect 4816 4137 4844 4168
rect 5000 4168 6929 4196
rect 4801 4131 4859 4137
rect 4801 4097 4813 4131
rect 4847 4097 4859 4131
rect 4801 4091 4859 4097
rect 4893 4131 4951 4137
rect 4893 4097 4905 4131
rect 4939 4128 4951 4131
rect 5000 4128 5028 4168
rect 6917 4165 6929 4168
rect 6963 4165 6975 4199
rect 6917 4159 6975 4165
rect 4939 4100 5028 4128
rect 5077 4131 5135 4137
rect 4939 4097 4951 4100
rect 4893 4091 4951 4097
rect 5077 4097 5089 4131
rect 5123 4128 5135 4131
rect 5258 4128 5264 4140
rect 5123 4100 5264 4128
rect 5123 4097 5135 4100
rect 5077 4091 5135 4097
rect 5258 4088 5264 4100
rect 5316 4088 5322 4140
rect 5350 4088 5356 4140
rect 5408 4088 5414 4140
rect 5445 4131 5503 4137
rect 5445 4097 5457 4131
rect 5491 4128 5503 4131
rect 5534 4128 5540 4140
rect 5491 4100 5540 4128
rect 5491 4097 5503 4100
rect 5445 4091 5503 4097
rect 5534 4088 5540 4100
rect 5592 4088 5598 4140
rect 5626 4088 5632 4140
rect 5684 4088 5690 4140
rect 6733 4131 6791 4137
rect 6733 4128 6745 4131
rect 5736 4100 6745 4128
rect 1504 4032 1900 4060
rect 2225 4063 2283 4069
rect 2225 4029 2237 4063
rect 2271 4060 2283 4063
rect 3789 4063 3847 4069
rect 3789 4060 3801 4063
rect 2271 4032 3801 4060
rect 2271 4029 2283 4032
rect 2225 4023 2283 4029
rect 3789 4029 3801 4032
rect 3835 4029 3847 4063
rect 5736 4060 5764 4100
rect 6733 4097 6745 4100
rect 6779 4128 6791 4131
rect 6822 4128 6828 4140
rect 6779 4100 6828 4128
rect 6779 4097 6791 4100
rect 6733 4091 6791 4097
rect 6822 4088 6828 4100
rect 6880 4088 6886 4140
rect 7193 4131 7251 4137
rect 7193 4128 7205 4131
rect 6932 4100 7205 4128
rect 3789 4023 3847 4029
rect 5276 4032 5764 4060
rect 3326 3952 3332 4004
rect 3384 3992 3390 4004
rect 3697 3995 3755 4001
rect 3697 3992 3709 3995
rect 3384 3964 3709 3992
rect 3384 3952 3390 3964
rect 3697 3961 3709 3964
rect 3743 3961 3755 3995
rect 3697 3955 3755 3961
rect 1857 3927 1915 3933
rect 1857 3893 1869 3927
rect 1903 3924 1915 3927
rect 2958 3924 2964 3936
rect 1903 3896 2964 3924
rect 1903 3893 1915 3896
rect 1857 3887 1915 3893
rect 2958 3884 2964 3896
rect 3016 3884 3022 3936
rect 3712 3924 3740 3955
rect 3970 3952 3976 4004
rect 4028 3992 4034 4004
rect 4065 3995 4123 4001
rect 4065 3992 4077 3995
rect 4028 3964 4077 3992
rect 4028 3952 4034 3964
rect 4065 3961 4077 3964
rect 4111 3961 4123 3995
rect 4065 3955 4123 3961
rect 4154 3952 4160 4004
rect 4212 3952 4218 4004
rect 4890 3952 4896 4004
rect 4948 3992 4954 4004
rect 4985 3995 5043 4001
rect 4985 3992 4997 3995
rect 4948 3964 4997 3992
rect 4948 3952 4954 3964
rect 4985 3961 4997 3964
rect 5031 3961 5043 3995
rect 4985 3955 5043 3961
rect 5276 3924 5304 4032
rect 6546 4020 6552 4072
rect 6604 4020 6610 4072
rect 6638 4020 6644 4072
rect 6696 4060 6702 4072
rect 6932 4060 6960 4100
rect 7193 4097 7205 4100
rect 7239 4097 7251 4131
rect 7193 4091 7251 4097
rect 6696 4032 6960 4060
rect 7101 4063 7159 4069
rect 6696 4020 6702 4032
rect 7101 4029 7113 4063
rect 7147 4029 7159 4063
rect 7101 4023 7159 4029
rect 7285 4063 7343 4069
rect 7285 4029 7297 4063
rect 7331 4029 7343 4063
rect 7285 4023 7343 4029
rect 5537 3995 5595 4001
rect 5537 3961 5549 3995
rect 5583 3992 5595 3995
rect 6365 3995 6423 4001
rect 6365 3992 6377 3995
rect 5583 3964 6377 3992
rect 5583 3961 5595 3964
rect 5537 3955 5595 3961
rect 6365 3961 6377 3964
rect 6411 3961 6423 3995
rect 6564 3992 6592 4020
rect 7116 3992 7144 4023
rect 6564 3964 7144 3992
rect 6365 3955 6423 3961
rect 7300 3936 7328 4023
rect 3712 3896 5304 3924
rect 5718 3884 5724 3936
rect 5776 3924 5782 3936
rect 5813 3927 5871 3933
rect 5813 3924 5825 3927
rect 5776 3896 5825 3924
rect 5776 3884 5782 3896
rect 5813 3893 5825 3896
rect 5859 3893 5871 3927
rect 5813 3887 5871 3893
rect 7282 3884 7288 3936
rect 7340 3884 7346 3936
rect 1104 3834 7912 3856
rect 1104 3782 1801 3834
rect 1853 3782 1865 3834
rect 1917 3782 1929 3834
rect 1981 3782 1993 3834
rect 2045 3782 2057 3834
rect 2109 3782 3503 3834
rect 3555 3782 3567 3834
rect 3619 3782 3631 3834
rect 3683 3782 3695 3834
rect 3747 3782 3759 3834
rect 3811 3782 5205 3834
rect 5257 3782 5269 3834
rect 5321 3782 5333 3834
rect 5385 3782 5397 3834
rect 5449 3782 5461 3834
rect 5513 3782 6907 3834
rect 6959 3782 6971 3834
rect 7023 3782 7035 3834
rect 7087 3782 7099 3834
rect 7151 3782 7163 3834
rect 7215 3782 7912 3834
rect 1104 3760 7912 3782
rect 2222 3720 2228 3732
rect 1780 3692 2228 3720
rect 1780 3593 1808 3692
rect 2222 3680 2228 3692
rect 2280 3680 2286 3732
rect 4154 3680 4160 3732
rect 4212 3680 4218 3732
rect 4706 3680 4712 3732
rect 4764 3680 4770 3732
rect 4985 3723 5043 3729
rect 4985 3689 4997 3723
rect 5031 3689 5043 3723
rect 4985 3683 5043 3689
rect 5261 3723 5319 3729
rect 5261 3689 5273 3723
rect 5307 3720 5319 3723
rect 5350 3720 5356 3732
rect 5307 3692 5356 3720
rect 5307 3689 5319 3692
rect 5261 3683 5319 3689
rect 4724 3652 4752 3680
rect 5000 3652 5028 3683
rect 5350 3680 5356 3692
rect 5408 3680 5414 3732
rect 4724 3624 5028 3652
rect 1765 3587 1823 3593
rect 1765 3553 1777 3587
rect 1811 3553 1823 3587
rect 1765 3547 1823 3553
rect 4798 3544 4804 3596
rect 4856 3584 4862 3596
rect 4985 3587 5043 3593
rect 4985 3584 4997 3587
rect 4856 3556 4997 3584
rect 4856 3544 4862 3556
rect 4985 3553 4997 3556
rect 5031 3553 5043 3587
rect 5353 3587 5411 3593
rect 5353 3584 5365 3587
rect 4985 3547 5043 3553
rect 5276 3556 5365 3584
rect 4062 3516 4068 3528
rect 3174 3488 4068 3516
rect 4062 3476 4068 3488
rect 4120 3476 4126 3528
rect 4341 3519 4399 3525
rect 4341 3485 4353 3519
rect 4387 3485 4399 3519
rect 4341 3479 4399 3485
rect 2041 3451 2099 3457
rect 2041 3417 2053 3451
rect 2087 3417 2099 3451
rect 2041 3411 2099 3417
rect 2056 3380 2084 3411
rect 3050 3380 3056 3392
rect 2056 3352 3056 3380
rect 3050 3340 3056 3352
rect 3108 3340 3114 3392
rect 3510 3340 3516 3392
rect 3568 3340 3574 3392
rect 4356 3380 4384 3479
rect 4522 3476 4528 3528
rect 4580 3476 4586 3528
rect 4617 3519 4675 3525
rect 4617 3485 4629 3519
rect 4663 3516 4675 3519
rect 4816 3516 4844 3544
rect 5276 3528 5304 3556
rect 5353 3553 5365 3556
rect 5399 3553 5411 3587
rect 5353 3547 5411 3553
rect 5629 3587 5687 3593
rect 5629 3553 5641 3587
rect 5675 3584 5687 3587
rect 5718 3584 5724 3596
rect 5675 3556 5724 3584
rect 5675 3553 5687 3556
rect 5629 3547 5687 3553
rect 5718 3544 5724 3556
rect 5776 3544 5782 3596
rect 4663 3488 4844 3516
rect 4916 3513 4974 3519
rect 4663 3485 4675 3488
rect 4617 3479 4675 3485
rect 4916 3479 4928 3513
rect 4962 3510 4974 3513
rect 4962 3482 5212 3510
rect 4962 3479 4974 3482
rect 4916 3473 4974 3479
rect 5184 3448 5212 3482
rect 5258 3476 5264 3528
rect 5316 3476 5322 3528
rect 7282 3516 7288 3528
rect 7116 3488 7288 3516
rect 5626 3448 5632 3460
rect 5184 3420 5632 3448
rect 5626 3408 5632 3420
rect 5684 3408 5690 3460
rect 6270 3408 6276 3460
rect 6328 3408 6334 3460
rect 6914 3380 6920 3392
rect 4356 3352 6920 3380
rect 6914 3340 6920 3352
rect 6972 3380 6978 3392
rect 7116 3389 7144 3488
rect 7282 3476 7288 3488
rect 7340 3476 7346 3528
rect 7101 3383 7159 3389
rect 7101 3380 7113 3383
rect 6972 3352 7113 3380
rect 6972 3340 6978 3352
rect 7101 3349 7113 3352
rect 7147 3349 7159 3383
rect 7101 3343 7159 3349
rect 7469 3383 7527 3389
rect 7469 3349 7481 3383
rect 7515 3380 7527 3383
rect 8018 3380 8024 3392
rect 7515 3352 8024 3380
rect 7515 3349 7527 3352
rect 7469 3343 7527 3349
rect 8018 3340 8024 3352
rect 8076 3340 8082 3392
rect 1104 3290 7912 3312
rect 1104 3238 2461 3290
rect 2513 3238 2525 3290
rect 2577 3238 2589 3290
rect 2641 3238 2653 3290
rect 2705 3238 2717 3290
rect 2769 3238 4163 3290
rect 4215 3238 4227 3290
rect 4279 3238 4291 3290
rect 4343 3238 4355 3290
rect 4407 3238 4419 3290
rect 4471 3238 5865 3290
rect 5917 3238 5929 3290
rect 5981 3238 5993 3290
rect 6045 3238 6057 3290
rect 6109 3238 6121 3290
rect 6173 3238 7567 3290
rect 7619 3238 7631 3290
rect 7683 3238 7695 3290
rect 7747 3238 7759 3290
rect 7811 3238 7823 3290
rect 7875 3238 7912 3290
rect 1104 3216 7912 3238
rect 4890 3136 4896 3188
rect 4948 3176 4954 3188
rect 5537 3179 5595 3185
rect 5537 3176 5549 3179
rect 4948 3148 5549 3176
rect 4948 3136 4954 3148
rect 5537 3145 5549 3148
rect 5583 3145 5595 3179
rect 5537 3139 5595 3145
rect 5626 3136 5632 3188
rect 5684 3176 5690 3188
rect 6365 3179 6423 3185
rect 6365 3176 6377 3179
rect 5684 3148 6377 3176
rect 5684 3136 5690 3148
rect 6365 3145 6377 3148
rect 6411 3145 6423 3179
rect 6365 3139 6423 3145
rect 6914 3136 6920 3188
rect 6972 3136 6978 3188
rect 4525 3111 4583 3117
rect 4525 3077 4537 3111
rect 4571 3108 4583 3111
rect 4982 3108 4988 3120
rect 4571 3080 4988 3108
rect 4571 3077 4583 3080
rect 4525 3071 4583 3077
rect 4982 3068 4988 3080
rect 5040 3068 5046 3120
rect 1397 3043 1455 3049
rect 1397 3040 1409 3043
rect 308 3012 1409 3040
rect 1397 3009 1409 3012
rect 1443 3009 1455 3043
rect 1397 3003 1455 3009
rect 3510 3000 3516 3052
rect 3568 3040 3574 3052
rect 5721 3043 5779 3049
rect 5721 3040 5733 3043
rect 3568 3012 5733 3040
rect 3568 3000 3574 3012
rect 5721 3009 5733 3012
rect 5767 3040 5779 3043
rect 5997 3043 6055 3049
rect 5767 3012 5856 3040
rect 5767 3009 5779 3012
rect 5721 3003 5779 3009
rect 1673 2975 1731 2981
rect 1673 2941 1685 2975
rect 1719 2972 1731 2975
rect 4522 2972 4528 2984
rect 1719 2944 4528 2972
rect 1719 2941 1731 2944
rect 1673 2935 1731 2941
rect 4522 2932 4528 2944
rect 4580 2932 4586 2984
rect 5074 2932 5080 2984
rect 5132 2932 5138 2984
rect 2314 2864 2320 2916
rect 2372 2904 2378 2916
rect 3237 2907 3295 2913
rect 3237 2904 3249 2907
rect 2372 2876 3249 2904
rect 2372 2864 2378 2876
rect 3237 2873 3249 2876
rect 3283 2904 3295 2907
rect 5092 2904 5120 2932
rect 3283 2876 5120 2904
rect 5828 2904 5856 3012
rect 5997 3009 6009 3043
rect 6043 3040 6055 3043
rect 6638 3040 6644 3052
rect 6043 3012 6644 3040
rect 6043 3009 6055 3012
rect 5997 3003 6055 3009
rect 6638 3000 6644 3012
rect 6696 3000 6702 3052
rect 6932 3049 6960 3136
rect 6917 3043 6975 3049
rect 6917 3009 6929 3043
rect 6963 3009 6975 3043
rect 6917 3003 6975 3009
rect 7285 3043 7343 3049
rect 7285 3009 7297 3043
rect 7331 3040 7343 3043
rect 7374 3040 7380 3052
rect 7331 3012 7380 3040
rect 7331 3009 7343 3012
rect 7285 3003 7343 3009
rect 7374 3000 7380 3012
rect 7432 3000 7438 3052
rect 5905 2975 5963 2981
rect 5905 2941 5917 2975
rect 5951 2972 5963 2975
rect 6546 2972 6552 2984
rect 5951 2944 6552 2972
rect 5951 2941 5963 2944
rect 5905 2935 5963 2941
rect 6546 2932 6552 2944
rect 6604 2932 6610 2984
rect 7282 2904 7288 2916
rect 5828 2876 7288 2904
rect 3283 2873 3295 2876
rect 3237 2867 3295 2873
rect 7282 2864 7288 2876
rect 7340 2864 7346 2916
rect 7469 2839 7527 2845
rect 7469 2805 7481 2839
rect 7515 2836 7527 2839
rect 8018 2836 8024 2848
rect 7515 2808 8024 2836
rect 7515 2805 7527 2808
rect 7469 2799 7527 2805
rect 8018 2796 8024 2808
rect 8076 2796 8082 2848
rect 1104 2746 7912 2768
rect 1104 2694 1801 2746
rect 1853 2694 1865 2746
rect 1917 2694 1929 2746
rect 1981 2694 1993 2746
rect 2045 2694 2057 2746
rect 2109 2694 3503 2746
rect 3555 2694 3567 2746
rect 3619 2694 3631 2746
rect 3683 2694 3695 2746
rect 3747 2694 3759 2746
rect 3811 2694 5205 2746
rect 5257 2694 5269 2746
rect 5321 2694 5333 2746
rect 5385 2694 5397 2746
rect 5449 2694 5461 2746
rect 5513 2694 6907 2746
rect 6959 2694 6971 2746
rect 7023 2694 7035 2746
rect 7087 2694 7099 2746
rect 7151 2694 7163 2746
rect 7215 2694 7912 2746
rect 1104 2672 7912 2694
rect 3973 2635 4031 2641
rect 3973 2601 3985 2635
rect 4019 2601 4031 2635
rect 3973 2595 4031 2601
rect 4157 2635 4215 2641
rect 4157 2601 4169 2635
rect 4203 2632 4215 2635
rect 4614 2632 4620 2644
rect 4203 2604 4620 2632
rect 4203 2601 4215 2604
rect 4157 2595 4215 2601
rect 3988 2564 4016 2595
rect 4614 2592 4620 2604
rect 4672 2592 4678 2644
rect 4706 2592 4712 2644
rect 4764 2592 4770 2644
rect 4724 2564 4752 2592
rect 3988 2536 4752 2564
rect 3326 2388 3332 2440
rect 3384 2428 3390 2440
rect 3789 2431 3847 2437
rect 3789 2428 3801 2431
rect 3384 2400 3801 2428
rect 3384 2388 3390 2400
rect 3789 2397 3801 2400
rect 3835 2397 3847 2431
rect 3789 2391 3847 2397
rect 3973 2431 4031 2437
rect 3973 2397 3985 2431
rect 4019 2428 4031 2431
rect 4798 2428 4804 2440
rect 4019 2400 4804 2428
rect 4019 2397 4031 2400
rect 3973 2391 4031 2397
rect 4798 2388 4804 2400
rect 4856 2388 4862 2440
rect 7009 2431 7067 2437
rect 7009 2397 7021 2431
rect 7055 2428 7067 2431
rect 7282 2428 7288 2440
rect 7055 2400 7288 2428
rect 7055 2397 7067 2400
rect 7009 2391 7067 2397
rect 7282 2388 7288 2400
rect 7340 2388 7346 2440
rect 6822 2252 6828 2304
rect 6880 2292 6886 2304
rect 7101 2295 7159 2301
rect 7101 2292 7113 2295
rect 6880 2264 7113 2292
rect 6880 2252 6886 2264
rect 7101 2261 7113 2264
rect 7147 2261 7159 2295
rect 7101 2255 7159 2261
rect 1104 2202 7912 2224
rect 1104 2150 2461 2202
rect 2513 2150 2525 2202
rect 2577 2150 2589 2202
rect 2641 2150 2653 2202
rect 2705 2150 2717 2202
rect 2769 2150 4163 2202
rect 4215 2150 4227 2202
rect 4279 2150 4291 2202
rect 4343 2150 4355 2202
rect 4407 2150 4419 2202
rect 4471 2150 5865 2202
rect 5917 2150 5929 2202
rect 5981 2150 5993 2202
rect 6045 2150 6057 2202
rect 6109 2150 6121 2202
rect 6173 2150 7567 2202
rect 7619 2150 7631 2202
rect 7683 2150 7695 2202
rect 7747 2150 7759 2202
rect 7811 2150 7823 2202
rect 7875 2150 7912 2202
rect 1104 2128 7912 2150
rect 388 1694 2934 1722
rect 388 1532 1804 1694
rect 2874 1532 2934 1694
rect 388 1512 2934 1532
rect 1764 1504 2934 1512
<< via1 >>
rect 2461 8678 2513 8730
rect 2525 8678 2577 8730
rect 2589 8678 2641 8730
rect 2653 8678 2705 8730
rect 2717 8678 2769 8730
rect 4163 8678 4215 8730
rect 4227 8678 4279 8730
rect 4291 8678 4343 8730
rect 4355 8678 4407 8730
rect 4419 8678 4471 8730
rect 5865 8678 5917 8730
rect 5929 8678 5981 8730
rect 5993 8678 6045 8730
rect 6057 8678 6109 8730
rect 6121 8678 6173 8730
rect 7567 8678 7619 8730
rect 7631 8678 7683 8730
rect 7695 8678 7747 8730
rect 7759 8678 7811 8730
rect 7823 8678 7875 8730
rect 6644 8619 6696 8628
rect 6644 8585 6653 8619
rect 6653 8585 6687 8619
rect 6687 8585 6696 8619
rect 6644 8576 6696 8585
rect 5080 8440 5132 8492
rect 7380 8440 7432 8492
rect 7472 8415 7524 8424
rect 7472 8381 7481 8415
rect 7481 8381 7515 8415
rect 7515 8381 7524 8415
rect 7472 8372 7524 8381
rect 2872 8304 2924 8356
rect 7288 8304 7340 8356
rect 2320 8279 2372 8288
rect 2320 8245 2329 8279
rect 2329 8245 2363 8279
rect 2363 8245 2372 8279
rect 2320 8236 2372 8245
rect 1801 8134 1853 8186
rect 1865 8134 1917 8186
rect 1929 8134 1981 8186
rect 1993 8134 2045 8186
rect 2057 8134 2109 8186
rect 3503 8134 3555 8186
rect 3567 8134 3619 8186
rect 3631 8134 3683 8186
rect 3695 8134 3747 8186
rect 3759 8134 3811 8186
rect 5205 8134 5257 8186
rect 5269 8134 5321 8186
rect 5333 8134 5385 8186
rect 5397 8134 5449 8186
rect 5461 8134 5513 8186
rect 6907 8134 6959 8186
rect 6971 8134 7023 8186
rect 7035 8134 7087 8186
rect 7099 8134 7151 8186
rect 7163 8134 7215 8186
rect 2320 8032 2372 8084
rect 6828 8032 6880 8084
rect 5540 7896 5592 7948
rect 2228 7760 2280 7812
rect 2872 7871 2924 7880
rect 2872 7837 2881 7871
rect 2881 7837 2915 7871
rect 2915 7837 2924 7871
rect 2872 7828 2924 7837
rect 4528 7871 4580 7880
rect 4528 7837 4537 7871
rect 4537 7837 4571 7871
rect 4571 7837 4580 7871
rect 4528 7828 4580 7837
rect 4896 7871 4948 7880
rect 4896 7837 4905 7871
rect 4905 7837 4939 7871
rect 4939 7837 4948 7871
rect 4896 7828 4948 7837
rect 1584 7735 1636 7744
rect 1584 7701 1593 7735
rect 1593 7701 1627 7735
rect 1627 7701 1636 7735
rect 1584 7692 1636 7701
rect 2964 7735 3016 7744
rect 2964 7701 2973 7735
rect 2973 7701 3007 7735
rect 3007 7701 3016 7735
rect 2964 7692 3016 7701
rect 4620 7692 4672 7744
rect 5264 7760 5316 7812
rect 6276 7760 6328 7812
rect 5724 7692 5776 7744
rect 6920 7692 6972 7744
rect 7472 7828 7524 7880
rect 8024 7692 8076 7744
rect 2461 7590 2513 7642
rect 2525 7590 2577 7642
rect 2589 7590 2641 7642
rect 2653 7590 2705 7642
rect 2717 7590 2769 7642
rect 4163 7590 4215 7642
rect 4227 7590 4279 7642
rect 4291 7590 4343 7642
rect 4355 7590 4407 7642
rect 4419 7590 4471 7642
rect 5865 7590 5917 7642
rect 5929 7590 5981 7642
rect 5993 7590 6045 7642
rect 6057 7590 6109 7642
rect 6121 7590 6173 7642
rect 7567 7590 7619 7642
rect 7631 7590 7683 7642
rect 7695 7590 7747 7642
rect 7759 7590 7811 7642
rect 7823 7590 7875 7642
rect 1584 7488 1636 7540
rect 6276 7488 6328 7540
rect 7932 7488 7984 7540
rect 4988 7463 5040 7472
rect 4988 7429 4997 7463
rect 4997 7429 5031 7463
rect 5031 7429 5040 7463
rect 4988 7420 5040 7429
rect 2320 7395 2372 7404
rect 2320 7361 2329 7395
rect 2329 7361 2363 7395
rect 2363 7361 2372 7395
rect 2320 7352 2372 7361
rect 4436 7395 4488 7404
rect 4436 7361 4445 7395
rect 4445 7361 4479 7395
rect 4479 7361 4488 7395
rect 4436 7352 4488 7361
rect 6920 7420 6972 7472
rect 7472 7352 7524 7404
rect 3332 7284 3384 7336
rect 3608 7284 3660 7336
rect 3976 7148 4028 7200
rect 4160 7191 4212 7200
rect 4160 7157 4169 7191
rect 4169 7157 4203 7191
rect 4203 7157 4212 7191
rect 4160 7148 4212 7157
rect 4896 7284 4948 7336
rect 5264 7327 5316 7336
rect 5264 7293 5273 7327
rect 5273 7293 5307 7327
rect 5307 7293 5316 7327
rect 5264 7284 5316 7293
rect 6368 7284 6420 7336
rect 6644 7284 6696 7336
rect 6920 7327 6972 7336
rect 6920 7293 6929 7327
rect 6929 7293 6963 7327
rect 6963 7293 6972 7327
rect 6920 7284 6972 7293
rect 5632 7148 5684 7200
rect 5816 7148 5868 7200
rect 1801 7046 1853 7098
rect 1865 7046 1917 7098
rect 1929 7046 1981 7098
rect 1993 7046 2045 7098
rect 2057 7046 2109 7098
rect 3503 7046 3555 7098
rect 3567 7046 3619 7098
rect 3631 7046 3683 7098
rect 3695 7046 3747 7098
rect 3759 7046 3811 7098
rect 5205 7046 5257 7098
rect 5269 7046 5321 7098
rect 5333 7046 5385 7098
rect 5397 7046 5449 7098
rect 5461 7046 5513 7098
rect 6907 7046 6959 7098
rect 6971 7046 7023 7098
rect 7035 7046 7087 7098
rect 7099 7046 7151 7098
rect 7163 7046 7215 7098
rect 2320 6944 2372 6996
rect 3700 6944 3752 6996
rect 4620 6944 4672 6996
rect 5632 6944 5684 6996
rect 7472 6944 7524 6996
rect 4160 6876 4212 6928
rect 4988 6876 5040 6928
rect 1584 6740 1636 6792
rect 3884 6740 3936 6792
rect 5540 6851 5592 6860
rect 5540 6817 5549 6851
rect 5549 6817 5583 6851
rect 5583 6817 5592 6851
rect 5540 6808 5592 6817
rect 5816 6808 5868 6860
rect 3056 6715 3108 6724
rect 3056 6681 3065 6715
rect 3065 6681 3099 6715
rect 3099 6681 3108 6715
rect 3056 6672 3108 6681
rect 3332 6672 3384 6724
rect 4068 6672 4120 6724
rect 1584 6647 1636 6656
rect 1584 6613 1593 6647
rect 1593 6613 1627 6647
rect 1627 6613 1636 6647
rect 1584 6604 1636 6613
rect 2872 6604 2924 6656
rect 3700 6604 3752 6656
rect 4528 6783 4580 6792
rect 4528 6749 4537 6783
rect 4537 6749 4571 6783
rect 4571 6749 4580 6783
rect 4528 6740 4580 6749
rect 4528 6604 4580 6656
rect 5172 6740 5224 6792
rect 5724 6672 5776 6724
rect 6276 6672 6328 6724
rect 4896 6604 4948 6656
rect 7380 6647 7432 6656
rect 7380 6613 7389 6647
rect 7389 6613 7423 6647
rect 7423 6613 7432 6647
rect 7380 6604 7432 6613
rect 2461 6502 2513 6554
rect 2525 6502 2577 6554
rect 2589 6502 2641 6554
rect 2653 6502 2705 6554
rect 2717 6502 2769 6554
rect 4163 6502 4215 6554
rect 4227 6502 4279 6554
rect 4291 6502 4343 6554
rect 4355 6502 4407 6554
rect 4419 6502 4471 6554
rect 5865 6502 5917 6554
rect 5929 6502 5981 6554
rect 5993 6502 6045 6554
rect 6057 6502 6109 6554
rect 6121 6502 6173 6554
rect 7567 6502 7619 6554
rect 7631 6502 7683 6554
rect 7695 6502 7747 6554
rect 7759 6502 7811 6554
rect 7823 6502 7875 6554
rect 3056 6400 3108 6452
rect 4068 6400 4120 6452
rect 5172 6400 5224 6452
rect 6368 6443 6420 6452
rect 6368 6409 6377 6443
rect 6377 6409 6411 6443
rect 6411 6409 6420 6443
rect 6368 6400 6420 6409
rect 2228 6264 2280 6316
rect 2596 6307 2648 6316
rect 2596 6273 2605 6307
rect 2605 6273 2639 6307
rect 2639 6273 2648 6307
rect 2596 6264 2648 6273
rect 2964 6332 3016 6384
rect 3884 6332 3936 6384
rect 4896 6332 4948 6384
rect 3148 6307 3200 6316
rect 3148 6273 3157 6307
rect 3157 6273 3191 6307
rect 3191 6273 3200 6307
rect 3148 6264 3200 6273
rect 4252 6264 4304 6316
rect 3516 6196 3568 6248
rect 3056 6171 3108 6180
rect 3056 6137 3065 6171
rect 3065 6137 3099 6171
rect 3099 6137 3108 6171
rect 3056 6128 3108 6137
rect 3976 6196 4028 6248
rect 6644 6332 6696 6384
rect 7104 6332 7156 6384
rect 6920 6264 6972 6316
rect 8024 6400 8076 6452
rect 7472 6264 7524 6316
rect 4804 6239 4856 6248
rect 3884 6128 3936 6180
rect 4804 6205 4813 6239
rect 4813 6205 4847 6239
rect 4847 6205 4856 6239
rect 4804 6196 4856 6205
rect 4896 6196 4948 6248
rect 2320 6060 2372 6112
rect 4344 6103 4396 6112
rect 4344 6069 4353 6103
rect 4353 6069 4387 6103
rect 4387 6069 4396 6103
rect 4344 6060 4396 6069
rect 1801 5958 1853 6010
rect 1865 5958 1917 6010
rect 1929 5958 1981 6010
rect 1993 5958 2045 6010
rect 2057 5958 2109 6010
rect 3503 5958 3555 6010
rect 3567 5958 3619 6010
rect 3631 5958 3683 6010
rect 3695 5958 3747 6010
rect 3759 5958 3811 6010
rect 5205 5958 5257 6010
rect 5269 5958 5321 6010
rect 5333 5958 5385 6010
rect 5397 5958 5449 6010
rect 5461 5958 5513 6010
rect 6907 5958 6959 6010
rect 6971 5958 7023 6010
rect 7035 5958 7087 6010
rect 7099 5958 7151 6010
rect 7163 5958 7215 6010
rect 2228 5856 2280 5908
rect 2872 5899 2924 5908
rect 2872 5865 2881 5899
rect 2881 5865 2915 5899
rect 2915 5865 2924 5899
rect 2872 5856 2924 5865
rect 3056 5856 3108 5908
rect 5080 5899 5132 5908
rect 5080 5865 5089 5899
rect 5089 5865 5123 5899
rect 5123 5865 5132 5899
rect 5080 5856 5132 5865
rect 4344 5788 4396 5840
rect 2596 5720 2648 5772
rect 4712 5720 4764 5772
rect 1584 5652 1636 5704
rect 3332 5695 3384 5704
rect 3332 5661 3341 5695
rect 3341 5661 3375 5695
rect 3375 5661 3384 5695
rect 3332 5652 3384 5661
rect 3516 5652 3568 5704
rect 3700 5652 3752 5704
rect 4252 5652 4304 5704
rect 2872 5584 2924 5636
rect 2964 5516 3016 5568
rect 3148 5516 3200 5568
rect 8024 5516 8076 5568
rect 2461 5414 2513 5466
rect 2525 5414 2577 5466
rect 2589 5414 2641 5466
rect 2653 5414 2705 5466
rect 2717 5414 2769 5466
rect 4163 5414 4215 5466
rect 4227 5414 4279 5466
rect 4291 5414 4343 5466
rect 4355 5414 4407 5466
rect 4419 5414 4471 5466
rect 5865 5414 5917 5466
rect 5929 5414 5981 5466
rect 5993 5414 6045 5466
rect 6057 5414 6109 5466
rect 6121 5414 6173 5466
rect 7567 5414 7619 5466
rect 7631 5414 7683 5466
rect 7695 5414 7747 5466
rect 7759 5414 7811 5466
rect 7823 5414 7875 5466
rect 2320 5312 2372 5364
rect 3516 5312 3568 5364
rect 3700 5312 3752 5364
rect 4528 5312 4580 5364
rect 2964 5244 3016 5296
rect 4160 5244 4212 5296
rect 3884 5176 3936 5228
rect 4068 5219 4120 5228
rect 4068 5185 4077 5219
rect 4077 5185 4111 5219
rect 4111 5185 4120 5219
rect 4068 5176 4120 5185
rect 4620 5176 4672 5228
rect 4804 5176 4856 5228
rect 7380 5176 7432 5228
rect 3424 5108 3476 5160
rect 3976 5108 4028 5160
rect 6276 5108 6328 5160
rect 4436 5040 4488 5092
rect 1584 5015 1636 5024
rect 1584 4981 1593 5015
rect 1593 4981 1627 5015
rect 1627 4981 1636 5015
rect 1584 4972 1636 4981
rect 2228 4972 2280 5024
rect 4896 4972 4948 5024
rect 5540 4972 5592 5024
rect 6552 4972 6604 5024
rect 1801 4870 1853 4922
rect 1865 4870 1917 4922
rect 1929 4870 1981 4922
rect 1993 4870 2045 4922
rect 2057 4870 2109 4922
rect 3503 4870 3555 4922
rect 3567 4870 3619 4922
rect 3631 4870 3683 4922
rect 3695 4870 3747 4922
rect 3759 4870 3811 4922
rect 5205 4870 5257 4922
rect 5269 4870 5321 4922
rect 5333 4870 5385 4922
rect 5397 4870 5449 4922
rect 5461 4870 5513 4922
rect 6907 4870 6959 4922
rect 6971 4870 7023 4922
rect 7035 4870 7087 4922
rect 7099 4870 7151 4922
rect 7163 4870 7215 4922
rect 2228 4811 2280 4820
rect 2228 4777 2237 4811
rect 2237 4777 2271 4811
rect 2271 4777 2280 4811
rect 2228 4768 2280 4777
rect 4896 4811 4948 4820
rect 4896 4777 4905 4811
rect 4905 4777 4939 4811
rect 4939 4777 4948 4811
rect 4896 4768 4948 4777
rect 2320 4675 2372 4684
rect 2320 4641 2329 4675
rect 2329 4641 2363 4675
rect 2363 4641 2372 4675
rect 2320 4632 2372 4641
rect 2964 4700 3016 4752
rect 3424 4700 3476 4752
rect 4436 4700 4488 4752
rect 3148 4496 3200 4548
rect 3884 4564 3936 4616
rect 4804 4632 4856 4684
rect 6644 4632 6696 4684
rect 6828 4632 6880 4684
rect 4528 4564 4580 4616
rect 5080 4564 5132 4616
rect 3056 4428 3108 4480
rect 3976 4428 4028 4480
rect 4160 4428 4212 4480
rect 4436 4428 4488 4480
rect 4712 4428 4764 4480
rect 4896 4428 4948 4480
rect 5264 4471 5316 4480
rect 5264 4437 5273 4471
rect 5273 4437 5307 4471
rect 5307 4437 5316 4471
rect 5264 4428 5316 4437
rect 5632 4539 5684 4548
rect 5632 4505 5641 4539
rect 5641 4505 5675 4539
rect 5675 4505 5684 4539
rect 5632 4496 5684 4505
rect 6276 4496 6328 4548
rect 7380 4428 7432 4480
rect 8024 4428 8076 4480
rect 2461 4326 2513 4378
rect 2525 4326 2577 4378
rect 2589 4326 2641 4378
rect 2653 4326 2705 4378
rect 2717 4326 2769 4378
rect 4163 4326 4215 4378
rect 4227 4326 4279 4378
rect 4291 4326 4343 4378
rect 4355 4326 4407 4378
rect 4419 4326 4471 4378
rect 5865 4326 5917 4378
rect 5929 4326 5981 4378
rect 5993 4326 6045 4378
rect 6057 4326 6109 4378
rect 6121 4326 6173 4378
rect 7567 4326 7619 4378
rect 7631 4326 7683 4378
rect 7695 4326 7747 4378
rect 7759 4326 7811 4378
rect 7823 4326 7875 4378
rect 1584 4224 1636 4276
rect 2228 4224 2280 4276
rect 3148 4224 3200 4276
rect 2320 4156 2372 4208
rect 5632 4224 5684 4276
rect 3884 4088 3936 4140
rect 4436 4156 4488 4208
rect 4620 4088 4672 4140
rect 5264 4088 5316 4140
rect 5356 4131 5408 4140
rect 5356 4097 5365 4131
rect 5365 4097 5399 4131
rect 5399 4097 5408 4131
rect 5356 4088 5408 4097
rect 5540 4088 5592 4140
rect 5632 4131 5684 4140
rect 5632 4097 5641 4131
rect 5641 4097 5675 4131
rect 5675 4097 5684 4131
rect 5632 4088 5684 4097
rect 6828 4088 6880 4140
rect 3332 3952 3384 4004
rect 2964 3884 3016 3936
rect 3976 3952 4028 4004
rect 4160 3995 4212 4004
rect 4160 3961 4169 3995
rect 4169 3961 4203 3995
rect 4203 3961 4212 3995
rect 4160 3952 4212 3961
rect 4896 3952 4948 4004
rect 6552 4063 6604 4072
rect 6552 4029 6561 4063
rect 6561 4029 6595 4063
rect 6595 4029 6604 4063
rect 6552 4020 6604 4029
rect 6644 4063 6696 4072
rect 6644 4029 6653 4063
rect 6653 4029 6687 4063
rect 6687 4029 6696 4063
rect 6644 4020 6696 4029
rect 5724 3884 5776 3936
rect 7288 3884 7340 3936
rect 1801 3782 1853 3834
rect 1865 3782 1917 3834
rect 1929 3782 1981 3834
rect 1993 3782 2045 3834
rect 2057 3782 2109 3834
rect 3503 3782 3555 3834
rect 3567 3782 3619 3834
rect 3631 3782 3683 3834
rect 3695 3782 3747 3834
rect 3759 3782 3811 3834
rect 5205 3782 5257 3834
rect 5269 3782 5321 3834
rect 5333 3782 5385 3834
rect 5397 3782 5449 3834
rect 5461 3782 5513 3834
rect 6907 3782 6959 3834
rect 6971 3782 7023 3834
rect 7035 3782 7087 3834
rect 7099 3782 7151 3834
rect 7163 3782 7215 3834
rect 2228 3680 2280 3732
rect 4160 3723 4212 3732
rect 4160 3689 4169 3723
rect 4169 3689 4203 3723
rect 4203 3689 4212 3723
rect 4160 3680 4212 3689
rect 4712 3680 4764 3732
rect 5356 3680 5408 3732
rect 4804 3544 4856 3596
rect 4068 3476 4120 3528
rect 3056 3340 3108 3392
rect 3516 3383 3568 3392
rect 3516 3349 3525 3383
rect 3525 3349 3559 3383
rect 3559 3349 3568 3383
rect 3516 3340 3568 3349
rect 4528 3519 4580 3528
rect 4528 3485 4537 3519
rect 4537 3485 4571 3519
rect 4571 3485 4580 3519
rect 4528 3476 4580 3485
rect 5724 3544 5776 3596
rect 5264 3476 5316 3528
rect 7288 3519 7340 3528
rect 5632 3408 5684 3460
rect 6276 3408 6328 3460
rect 6920 3340 6972 3392
rect 7288 3485 7297 3519
rect 7297 3485 7331 3519
rect 7331 3485 7340 3519
rect 7288 3476 7340 3485
rect 8024 3340 8076 3392
rect 2461 3238 2513 3290
rect 2525 3238 2577 3290
rect 2589 3238 2641 3290
rect 2653 3238 2705 3290
rect 2717 3238 2769 3290
rect 4163 3238 4215 3290
rect 4227 3238 4279 3290
rect 4291 3238 4343 3290
rect 4355 3238 4407 3290
rect 4419 3238 4471 3290
rect 5865 3238 5917 3290
rect 5929 3238 5981 3290
rect 5993 3238 6045 3290
rect 6057 3238 6109 3290
rect 6121 3238 6173 3290
rect 7567 3238 7619 3290
rect 7631 3238 7683 3290
rect 7695 3238 7747 3290
rect 7759 3238 7811 3290
rect 7823 3238 7875 3290
rect 4896 3136 4948 3188
rect 5632 3136 5684 3188
rect 6920 3136 6972 3188
rect 4988 3068 5040 3120
rect 3516 3000 3568 3052
rect 4528 2932 4580 2984
rect 5080 2932 5132 2984
rect 2320 2864 2372 2916
rect 6644 3000 6696 3052
rect 7380 3000 7432 3052
rect 6552 2932 6604 2984
rect 7288 2864 7340 2916
rect 8024 2796 8076 2848
rect 1801 2694 1853 2746
rect 1865 2694 1917 2746
rect 1929 2694 1981 2746
rect 1993 2694 2045 2746
rect 2057 2694 2109 2746
rect 3503 2694 3555 2746
rect 3567 2694 3619 2746
rect 3631 2694 3683 2746
rect 3695 2694 3747 2746
rect 3759 2694 3811 2746
rect 5205 2694 5257 2746
rect 5269 2694 5321 2746
rect 5333 2694 5385 2746
rect 5397 2694 5449 2746
rect 5461 2694 5513 2746
rect 6907 2694 6959 2746
rect 6971 2694 7023 2746
rect 7035 2694 7087 2746
rect 7099 2694 7151 2746
rect 7163 2694 7215 2746
rect 4620 2592 4672 2644
rect 4712 2592 4764 2644
rect 3332 2388 3384 2440
rect 4804 2388 4856 2440
rect 7288 2388 7340 2440
rect 6828 2252 6880 2304
rect 2461 2150 2513 2202
rect 2525 2150 2577 2202
rect 2589 2150 2641 2202
rect 2653 2150 2705 2202
rect 2717 2150 2769 2202
rect 4163 2150 4215 2202
rect 4227 2150 4279 2202
rect 4291 2150 4343 2202
rect 4355 2150 4407 2202
rect 4419 2150 4471 2202
rect 5865 2150 5917 2202
rect 5929 2150 5981 2202
rect 5993 2150 6045 2202
rect 6057 2150 6109 2202
rect 6121 2150 6173 2202
rect 7567 2150 7619 2202
rect 7631 2150 7683 2202
rect 7695 2150 7747 2202
rect 7759 2150 7811 2202
rect 7823 2150 7875 2202
rect 1804 1532 2874 1694
<< metal2 >>
rect 6642 9888 6698 9897
rect 6642 9823 6698 9832
rect 2461 8732 2769 8741
rect 2461 8730 2467 8732
rect 2523 8730 2547 8732
rect 2603 8730 2627 8732
rect 2683 8730 2707 8732
rect 2763 8730 2769 8732
rect 2523 8678 2525 8730
rect 2705 8678 2707 8730
rect 2461 8676 2467 8678
rect 2523 8676 2547 8678
rect 2603 8676 2627 8678
rect 2683 8676 2707 8678
rect 2763 8676 2769 8678
rect 2461 8667 2769 8676
rect 4163 8732 4471 8741
rect 4163 8730 4169 8732
rect 4225 8730 4249 8732
rect 4305 8730 4329 8732
rect 4385 8730 4409 8732
rect 4465 8730 4471 8732
rect 4225 8678 4227 8730
rect 4407 8678 4409 8730
rect 4163 8676 4169 8678
rect 4225 8676 4249 8678
rect 4305 8676 4329 8678
rect 4385 8676 4409 8678
rect 4465 8676 4471 8678
rect 4163 8667 4471 8676
rect 5865 8732 6173 8741
rect 5865 8730 5871 8732
rect 5927 8730 5951 8732
rect 6007 8730 6031 8732
rect 6087 8730 6111 8732
rect 6167 8730 6173 8732
rect 5927 8678 5929 8730
rect 6109 8678 6111 8730
rect 5865 8676 5871 8678
rect 5927 8676 5951 8678
rect 6007 8676 6031 8678
rect 6087 8676 6111 8678
rect 6167 8676 6173 8678
rect 5865 8667 6173 8676
rect 6656 8634 6684 9823
rect 8022 8800 8078 8809
rect 7944 8758 8022 8786
rect 7567 8732 7875 8741
rect 7567 8730 7573 8732
rect 7629 8730 7653 8732
rect 7709 8730 7733 8732
rect 7789 8730 7813 8732
rect 7869 8730 7875 8732
rect 7629 8678 7631 8730
rect 7811 8678 7813 8730
rect 7567 8676 7573 8678
rect 7629 8676 7653 8678
rect 7709 8676 7733 8678
rect 7789 8676 7813 8678
rect 7869 8676 7875 8678
rect 7567 8667 7875 8676
rect 6644 8628 6696 8634
rect 6644 8570 6696 8576
rect 5080 8492 5132 8498
rect 5080 8434 5132 8440
rect 7380 8492 7432 8498
rect 7380 8434 7432 8440
rect 2872 8356 2924 8362
rect 2872 8298 2924 8304
rect 2320 8288 2372 8294
rect 2320 8230 2372 8236
rect 1801 8188 2109 8197
rect 1801 8186 1807 8188
rect 1863 8186 1887 8188
rect 1943 8186 1967 8188
rect 2023 8186 2047 8188
rect 2103 8186 2109 8188
rect 1863 8134 1865 8186
rect 2045 8134 2047 8186
rect 1801 8132 1807 8134
rect 1863 8132 1887 8134
rect 1943 8132 1967 8134
rect 2023 8132 2047 8134
rect 2103 8132 2109 8134
rect 1801 8123 2109 8132
rect 2332 8090 2360 8230
rect 2320 8084 2372 8090
rect 2320 8026 2372 8032
rect 2228 7812 2280 7818
rect 2228 7754 2280 7760
rect 1584 7744 1636 7750
rect 1584 7686 1636 7692
rect 1596 7546 1624 7686
rect 1584 7540 1636 7546
rect 1584 7482 1636 7488
rect 1596 6798 1624 7482
rect 1801 7100 2109 7109
rect 1801 7098 1807 7100
rect 1863 7098 1887 7100
rect 1943 7098 1967 7100
rect 2023 7098 2047 7100
rect 2103 7098 2109 7100
rect 1863 7046 1865 7098
rect 2045 7046 2047 7098
rect 1801 7044 1807 7046
rect 1863 7044 1887 7046
rect 1943 7044 1967 7046
rect 2023 7044 2047 7046
rect 2103 7044 2109 7046
rect 1801 7035 2109 7044
rect 1584 6792 1636 6798
rect 1584 6734 1636 6740
rect 1584 6656 1636 6662
rect 1584 6598 1636 6604
rect 1596 5710 1624 6598
rect 2240 6322 2268 7754
rect 2332 7410 2360 8026
rect 2884 7886 2912 8298
rect 3503 8188 3811 8197
rect 3503 8186 3509 8188
rect 3565 8186 3589 8188
rect 3645 8186 3669 8188
rect 3725 8186 3749 8188
rect 3805 8186 3811 8188
rect 3565 8134 3567 8186
rect 3747 8134 3749 8186
rect 3503 8132 3509 8134
rect 3565 8132 3589 8134
rect 3645 8132 3669 8134
rect 3725 8132 3749 8134
rect 3805 8132 3811 8134
rect 3503 8123 3811 8132
rect 2872 7880 2924 7886
rect 2872 7822 2924 7828
rect 4528 7880 4580 7886
rect 4528 7822 4580 7828
rect 4896 7880 4948 7886
rect 4896 7822 4948 7828
rect 2461 7644 2769 7653
rect 2461 7642 2467 7644
rect 2523 7642 2547 7644
rect 2603 7642 2627 7644
rect 2683 7642 2707 7644
rect 2763 7642 2769 7644
rect 2523 7590 2525 7642
rect 2705 7590 2707 7642
rect 2461 7588 2467 7590
rect 2523 7588 2547 7590
rect 2603 7588 2627 7590
rect 2683 7588 2707 7590
rect 2763 7588 2769 7590
rect 2461 7579 2769 7588
rect 2320 7404 2372 7410
rect 2320 7346 2372 7352
rect 2332 7002 2360 7346
rect 2320 6996 2372 7002
rect 2320 6938 2372 6944
rect 2884 6662 2912 7822
rect 2964 7744 3016 7750
rect 2964 7686 3016 7692
rect 2872 6656 2924 6662
rect 2872 6598 2924 6604
rect 2461 6556 2769 6565
rect 2461 6554 2467 6556
rect 2523 6554 2547 6556
rect 2603 6554 2627 6556
rect 2683 6554 2707 6556
rect 2763 6554 2769 6556
rect 2523 6502 2525 6554
rect 2705 6502 2707 6554
rect 2461 6500 2467 6502
rect 2523 6500 2547 6502
rect 2603 6500 2627 6502
rect 2683 6500 2707 6502
rect 2763 6500 2769 6502
rect 2461 6491 2769 6500
rect 2228 6316 2280 6322
rect 2228 6258 2280 6264
rect 2596 6316 2648 6322
rect 2596 6258 2648 6264
rect 2320 6112 2372 6118
rect 2320 6054 2372 6060
rect 1801 6012 2109 6021
rect 1801 6010 1807 6012
rect 1863 6010 1887 6012
rect 1943 6010 1967 6012
rect 2023 6010 2047 6012
rect 2103 6010 2109 6012
rect 1863 5958 1865 6010
rect 2045 5958 2047 6010
rect 1801 5956 1807 5958
rect 1863 5956 1887 5958
rect 1943 5956 1967 5958
rect 2023 5956 2047 5958
rect 2103 5956 2109 5958
rect 1801 5947 2109 5956
rect 2228 5908 2280 5914
rect 2228 5850 2280 5856
rect 1584 5704 1636 5710
rect 1584 5646 1636 5652
rect 2240 5030 2268 5850
rect 2332 5370 2360 6054
rect 2608 5778 2636 6258
rect 2884 5914 2912 6598
rect 2976 6390 3004 7686
rect 4163 7644 4471 7653
rect 4163 7642 4169 7644
rect 4225 7642 4249 7644
rect 4305 7642 4329 7644
rect 4385 7642 4409 7644
rect 4465 7642 4471 7644
rect 4225 7590 4227 7642
rect 4407 7590 4409 7642
rect 4163 7588 4169 7590
rect 4225 7588 4249 7590
rect 4305 7588 4329 7590
rect 4385 7588 4409 7590
rect 4465 7588 4471 7590
rect 4163 7579 4471 7588
rect 4434 7440 4490 7449
rect 4434 7375 4436 7384
rect 4488 7375 4490 7384
rect 4436 7346 4488 7352
rect 3332 7336 3384 7342
rect 3608 7336 3660 7342
rect 3332 7278 3384 7284
rect 3436 7296 3608 7324
rect 3344 6730 3372 7278
rect 3056 6724 3108 6730
rect 3056 6666 3108 6672
rect 3332 6724 3384 6730
rect 3332 6666 3384 6672
rect 3068 6458 3096 6666
rect 3056 6452 3108 6458
rect 3056 6394 3108 6400
rect 2964 6384 3016 6390
rect 2964 6326 3016 6332
rect 2872 5908 2924 5914
rect 2872 5850 2924 5856
rect 2596 5772 2648 5778
rect 2596 5714 2648 5720
rect 2976 5658 3004 6326
rect 3148 6316 3200 6322
rect 3148 6258 3200 6264
rect 3056 6180 3108 6186
rect 3056 6122 3108 6128
rect 3068 5914 3096 6122
rect 3056 5908 3108 5914
rect 3056 5850 3108 5856
rect 2872 5636 2924 5642
rect 2976 5630 3096 5658
rect 2872 5578 2924 5584
rect 2461 5468 2769 5477
rect 2461 5466 2467 5468
rect 2523 5466 2547 5468
rect 2603 5466 2627 5468
rect 2683 5466 2707 5468
rect 2763 5466 2769 5468
rect 2523 5414 2525 5466
rect 2705 5414 2707 5466
rect 2461 5412 2467 5414
rect 2523 5412 2547 5414
rect 2603 5412 2627 5414
rect 2683 5412 2707 5414
rect 2763 5412 2769 5414
rect 2461 5403 2769 5412
rect 2320 5364 2372 5370
rect 2320 5306 2372 5312
rect 1584 5024 1636 5030
rect 1584 4966 1636 4972
rect 2228 5024 2280 5030
rect 2228 4966 2280 4972
rect 1596 4282 1624 4966
rect 1801 4924 2109 4933
rect 1801 4922 1807 4924
rect 1863 4922 1887 4924
rect 1943 4922 1967 4924
rect 2023 4922 2047 4924
rect 2103 4922 2109 4924
rect 1863 4870 1865 4922
rect 2045 4870 2047 4922
rect 1801 4868 1807 4870
rect 1863 4868 1887 4870
rect 1943 4868 1967 4870
rect 2023 4868 2047 4870
rect 2103 4868 2109 4870
rect 1801 4859 2109 4868
rect 2240 4826 2268 4966
rect 2228 4820 2280 4826
rect 2228 4762 2280 4768
rect 2332 4690 2360 5306
rect 2320 4684 2372 4690
rect 2240 4644 2320 4672
rect 2240 4282 2268 4644
rect 2320 4626 2372 4632
rect 2461 4380 2769 4389
rect 2461 4378 2467 4380
rect 2523 4378 2547 4380
rect 2603 4378 2627 4380
rect 2683 4378 2707 4380
rect 2763 4378 2769 4380
rect 2523 4326 2525 4378
rect 2705 4326 2707 4378
rect 2461 4324 2467 4326
rect 2523 4324 2547 4326
rect 2603 4324 2627 4326
rect 2683 4324 2707 4326
rect 2763 4324 2769 4326
rect 2461 4315 2769 4324
rect 1584 4276 1636 4282
rect 1584 4218 1636 4224
rect 2228 4276 2280 4282
rect 2228 4218 2280 4224
rect 2320 4208 2372 4214
rect 2320 4150 2372 4156
rect 1801 3836 2109 3845
rect 1801 3834 1807 3836
rect 1863 3834 1887 3836
rect 1943 3834 1967 3836
rect 2023 3834 2047 3836
rect 2103 3834 2109 3836
rect 1863 3782 1865 3834
rect 2045 3782 2047 3834
rect 1801 3780 1807 3782
rect 1863 3780 1887 3782
rect 1943 3780 1967 3782
rect 2023 3780 2047 3782
rect 2103 3780 2109 3782
rect 1801 3771 2109 3780
rect 2228 3732 2280 3738
rect 2332 3720 2360 4150
rect 2280 3692 2360 3720
rect 2228 3674 2280 3680
rect 2332 2922 2360 3692
rect 2461 3292 2769 3301
rect 2461 3290 2467 3292
rect 2523 3290 2547 3292
rect 2603 3290 2627 3292
rect 2683 3290 2707 3292
rect 2763 3290 2769 3292
rect 2523 3238 2525 3290
rect 2705 3238 2707 3290
rect 2461 3236 2467 3238
rect 2523 3236 2547 3238
rect 2603 3236 2627 3238
rect 2683 3236 2707 3238
rect 2763 3236 2769 3238
rect 2461 3227 2769 3236
rect 2320 2916 2372 2922
rect 2320 2858 2372 2864
rect 1801 2748 2109 2757
rect 1801 2746 1807 2748
rect 1863 2746 1887 2748
rect 1943 2746 1967 2748
rect 2023 2746 2047 2748
rect 2103 2746 2109 2748
rect 1863 2694 1865 2746
rect 2045 2694 2047 2746
rect 1801 2692 1807 2694
rect 1863 2692 1887 2694
rect 1943 2692 1967 2694
rect 2023 2692 2047 2694
rect 2103 2692 2109 2694
rect 1801 2683 2109 2692
rect 2461 2204 2769 2213
rect 2461 2202 2467 2204
rect 2523 2202 2547 2204
rect 2603 2202 2627 2204
rect 2683 2202 2707 2204
rect 2763 2202 2769 2204
rect 2523 2150 2525 2202
rect 2705 2150 2707 2202
rect 2461 2148 2467 2150
rect 2523 2148 2547 2150
rect 2603 2148 2627 2150
rect 2683 2148 2707 2150
rect 2763 2148 2769 2150
rect 2461 2139 2769 2148
rect 2884 1718 2912 5578
rect 2964 5568 3016 5574
rect 2964 5510 3016 5516
rect 2976 5302 3004 5510
rect 2964 5296 3016 5302
rect 2964 5238 3016 5244
rect 2964 4752 3016 4758
rect 2964 4694 3016 4700
rect 2976 3942 3004 4694
rect 3068 4570 3096 5630
rect 3160 5574 3188 6258
rect 3436 6236 3464 7296
rect 3608 7278 3660 7284
rect 3976 7200 4028 7206
rect 3976 7142 4028 7148
rect 4160 7200 4212 7206
rect 4160 7142 4212 7148
rect 3503 7100 3811 7109
rect 3503 7098 3509 7100
rect 3565 7098 3589 7100
rect 3645 7098 3669 7100
rect 3725 7098 3749 7100
rect 3805 7098 3811 7100
rect 3565 7046 3567 7098
rect 3747 7046 3749 7098
rect 3503 7044 3509 7046
rect 3565 7044 3589 7046
rect 3645 7044 3669 7046
rect 3725 7044 3749 7046
rect 3805 7044 3811 7046
rect 3503 7035 3811 7044
rect 3700 6996 3752 7002
rect 3700 6938 3752 6944
rect 3712 6662 3740 6938
rect 3884 6792 3936 6798
rect 3884 6734 3936 6740
rect 3700 6656 3752 6662
rect 3700 6598 3752 6604
rect 3896 6390 3924 6734
rect 3884 6384 3936 6390
rect 3884 6326 3936 6332
rect 3988 6254 4016 7142
rect 4172 6934 4200 7142
rect 4160 6928 4212 6934
rect 4160 6870 4212 6876
rect 4540 6798 4568 7822
rect 4620 7744 4672 7750
rect 4620 7686 4672 7692
rect 4632 7002 4660 7686
rect 4908 7342 4936 7822
rect 4988 7472 5040 7478
rect 4988 7414 5040 7420
rect 4896 7336 4948 7342
rect 4896 7278 4948 7284
rect 4620 6996 4672 7002
rect 4620 6938 4672 6944
rect 5000 6934 5028 7414
rect 4988 6928 5040 6934
rect 4988 6870 5040 6876
rect 4528 6792 4580 6798
rect 4580 6740 4660 6746
rect 4528 6734 4660 6740
rect 4068 6724 4120 6730
rect 4540 6718 4660 6734
rect 4068 6666 4120 6672
rect 4080 6458 4108 6666
rect 4528 6656 4580 6662
rect 4528 6598 4580 6604
rect 4163 6556 4471 6565
rect 4163 6554 4169 6556
rect 4225 6554 4249 6556
rect 4305 6554 4329 6556
rect 4385 6554 4409 6556
rect 4465 6554 4471 6556
rect 4225 6502 4227 6554
rect 4407 6502 4409 6554
rect 4163 6500 4169 6502
rect 4225 6500 4249 6502
rect 4305 6500 4329 6502
rect 4385 6500 4409 6502
rect 4465 6500 4471 6502
rect 4163 6491 4471 6500
rect 4068 6452 4120 6458
rect 4068 6394 4120 6400
rect 4252 6316 4304 6322
rect 4252 6258 4304 6264
rect 3516 6248 3568 6254
rect 3436 6208 3516 6236
rect 3332 5704 3384 5710
rect 3332 5646 3384 5652
rect 3148 5568 3200 5574
rect 3148 5510 3200 5516
rect 3068 4554 3188 4570
rect 3068 4548 3200 4554
rect 3068 4542 3148 4548
rect 3148 4490 3200 4496
rect 3056 4480 3108 4486
rect 3056 4422 3108 4428
rect 2964 3936 3016 3942
rect 2964 3878 3016 3884
rect 3068 3398 3096 4422
rect 3160 4282 3188 4490
rect 3148 4276 3200 4282
rect 3148 4218 3200 4224
rect 3344 4010 3372 5646
rect 3436 5166 3464 6208
rect 3516 6190 3568 6196
rect 3976 6248 4028 6254
rect 3976 6190 4028 6196
rect 3884 6180 3936 6186
rect 3884 6122 3936 6128
rect 3503 6012 3811 6021
rect 3503 6010 3509 6012
rect 3565 6010 3589 6012
rect 3645 6010 3669 6012
rect 3725 6010 3749 6012
rect 3805 6010 3811 6012
rect 3565 5958 3567 6010
rect 3747 5958 3749 6010
rect 3503 5956 3509 5958
rect 3565 5956 3589 5958
rect 3645 5956 3669 5958
rect 3725 5956 3749 5958
rect 3805 5956 3811 5958
rect 3503 5947 3811 5956
rect 3516 5704 3568 5710
rect 3516 5646 3568 5652
rect 3700 5704 3752 5710
rect 3700 5646 3752 5652
rect 3528 5370 3556 5646
rect 3712 5370 3740 5646
rect 3516 5364 3568 5370
rect 3516 5306 3568 5312
rect 3700 5364 3752 5370
rect 3700 5306 3752 5312
rect 3896 5234 3924 6122
rect 3988 5556 4016 6190
rect 4264 5710 4292 6258
rect 4344 6112 4396 6118
rect 4344 6054 4396 6060
rect 4356 5846 4384 6054
rect 4344 5840 4396 5846
rect 4344 5782 4396 5788
rect 4252 5704 4304 5710
rect 4252 5646 4304 5652
rect 3988 5528 4108 5556
rect 4080 5234 4108 5528
rect 4163 5468 4471 5477
rect 4163 5466 4169 5468
rect 4225 5466 4249 5468
rect 4305 5466 4329 5468
rect 4385 5466 4409 5468
rect 4465 5466 4471 5468
rect 4225 5414 4227 5466
rect 4407 5414 4409 5466
rect 4163 5412 4169 5414
rect 4225 5412 4249 5414
rect 4305 5412 4329 5414
rect 4385 5412 4409 5414
rect 4465 5412 4471 5414
rect 4163 5403 4471 5412
rect 4540 5370 4568 6598
rect 4528 5364 4580 5370
rect 4528 5306 4580 5312
rect 4160 5296 4212 5302
rect 4160 5238 4212 5244
rect 3884 5228 3936 5234
rect 3884 5170 3936 5176
rect 4068 5228 4120 5234
rect 4068 5170 4120 5176
rect 3424 5160 3476 5166
rect 3424 5102 3476 5108
rect 3503 4924 3811 4933
rect 3503 4922 3509 4924
rect 3565 4922 3589 4924
rect 3645 4922 3669 4924
rect 3725 4922 3749 4924
rect 3805 4922 3811 4924
rect 3565 4870 3567 4922
rect 3747 4870 3749 4922
rect 3503 4868 3509 4870
rect 3565 4868 3589 4870
rect 3645 4868 3669 4870
rect 3725 4868 3749 4870
rect 3805 4868 3811 4870
rect 3503 4859 3811 4868
rect 3424 4752 3476 4758
rect 3424 4694 3476 4700
rect 3332 4004 3384 4010
rect 3332 3946 3384 3952
rect 3056 3392 3108 3398
rect 3056 3334 3108 3340
rect 3344 2446 3372 3946
rect 3436 3618 3464 4694
rect 3896 4622 3924 5170
rect 3976 5160 4028 5166
rect 4028 5108 4108 5114
rect 3976 5102 4108 5108
rect 3988 5086 4108 5102
rect 3884 4616 3936 4622
rect 3884 4558 3936 4564
rect 3976 4480 4028 4486
rect 3976 4422 4028 4428
rect 3884 4140 3936 4146
rect 3884 4082 3936 4088
rect 3896 3890 3924 4082
rect 3988 4010 4016 4422
rect 3976 4004 4028 4010
rect 3976 3946 4028 3952
rect 4080 3890 4108 5086
rect 4172 4486 4200 5238
rect 4632 5234 4660 6718
rect 4896 6656 4948 6662
rect 4896 6598 4948 6604
rect 4908 6390 4936 6598
rect 4896 6384 4948 6390
rect 4896 6326 4948 6332
rect 4804 6248 4856 6254
rect 4804 6190 4856 6196
rect 4896 6248 4948 6254
rect 4896 6190 4948 6196
rect 4712 5772 4764 5778
rect 4712 5714 4764 5720
rect 4620 5228 4672 5234
rect 4620 5170 4672 5176
rect 4436 5092 4488 5098
rect 4436 5034 4488 5040
rect 4448 4758 4476 5034
rect 4436 4752 4488 4758
rect 4436 4694 4488 4700
rect 4448 4486 4476 4694
rect 4528 4616 4580 4622
rect 4724 4604 4752 5714
rect 4816 5234 4844 6190
rect 4804 5228 4856 5234
rect 4804 5170 4856 5176
rect 4816 4690 4844 5170
rect 4908 5030 4936 6190
rect 5092 5914 5120 8434
rect 7288 8356 7340 8362
rect 7288 8298 7340 8304
rect 5205 8188 5513 8197
rect 5205 8186 5211 8188
rect 5267 8186 5291 8188
rect 5347 8186 5371 8188
rect 5427 8186 5451 8188
rect 5507 8186 5513 8188
rect 5267 8134 5269 8186
rect 5449 8134 5451 8186
rect 5205 8132 5211 8134
rect 5267 8132 5291 8134
rect 5347 8132 5371 8134
rect 5427 8132 5451 8134
rect 5507 8132 5513 8134
rect 5205 8123 5513 8132
rect 6907 8188 7215 8197
rect 6907 8186 6913 8188
rect 6969 8186 6993 8188
rect 7049 8186 7073 8188
rect 7129 8186 7153 8188
rect 7209 8186 7215 8188
rect 6969 8134 6971 8186
rect 7151 8134 7153 8186
rect 6907 8132 6913 8134
rect 6969 8132 6993 8134
rect 7049 8132 7073 8134
rect 7129 8132 7153 8134
rect 7209 8132 7215 8134
rect 6907 8123 7215 8132
rect 6828 8084 6880 8090
rect 6828 8026 6880 8032
rect 5540 7948 5592 7954
rect 5540 7890 5592 7896
rect 5264 7812 5316 7818
rect 5264 7754 5316 7760
rect 5276 7449 5304 7754
rect 5262 7440 5318 7449
rect 5262 7375 5318 7384
rect 5276 7342 5304 7375
rect 5264 7336 5316 7342
rect 5264 7278 5316 7284
rect 5205 7100 5513 7109
rect 5205 7098 5211 7100
rect 5267 7098 5291 7100
rect 5347 7098 5371 7100
rect 5427 7098 5451 7100
rect 5507 7098 5513 7100
rect 5267 7046 5269 7098
rect 5449 7046 5451 7098
rect 5205 7044 5211 7046
rect 5267 7044 5291 7046
rect 5347 7044 5371 7046
rect 5427 7044 5451 7046
rect 5507 7044 5513 7046
rect 5205 7035 5513 7044
rect 5552 6866 5580 7890
rect 6276 7812 6328 7818
rect 6276 7754 6328 7760
rect 5724 7744 5776 7750
rect 5724 7686 5776 7692
rect 5632 7200 5684 7206
rect 5632 7142 5684 7148
rect 5644 7002 5672 7142
rect 5632 6996 5684 7002
rect 5632 6938 5684 6944
rect 5540 6860 5592 6866
rect 5540 6802 5592 6808
rect 5172 6792 5224 6798
rect 5172 6734 5224 6740
rect 5184 6458 5212 6734
rect 5736 6730 5764 7686
rect 5865 7644 6173 7653
rect 5865 7642 5871 7644
rect 5927 7642 5951 7644
rect 6007 7642 6031 7644
rect 6087 7642 6111 7644
rect 6167 7642 6173 7644
rect 5927 7590 5929 7642
rect 6109 7590 6111 7642
rect 5865 7588 5871 7590
rect 5927 7588 5951 7590
rect 6007 7588 6031 7590
rect 6087 7588 6111 7590
rect 6167 7588 6173 7590
rect 5865 7579 6173 7588
rect 6288 7546 6316 7754
rect 6276 7540 6328 7546
rect 6276 7482 6328 7488
rect 5816 7200 5868 7206
rect 5816 7142 5868 7148
rect 5828 6866 5856 7142
rect 5816 6860 5868 6866
rect 5816 6802 5868 6808
rect 6288 6730 6316 7482
rect 6368 7336 6420 7342
rect 6368 7278 6420 7284
rect 6644 7336 6696 7342
rect 6644 7278 6696 7284
rect 5724 6724 5776 6730
rect 5724 6666 5776 6672
rect 6276 6724 6328 6730
rect 6276 6666 6328 6672
rect 5865 6556 6173 6565
rect 5865 6554 5871 6556
rect 5927 6554 5951 6556
rect 6007 6554 6031 6556
rect 6087 6554 6111 6556
rect 6167 6554 6173 6556
rect 5927 6502 5929 6554
rect 6109 6502 6111 6554
rect 5865 6500 5871 6502
rect 5927 6500 5951 6502
rect 6007 6500 6031 6502
rect 6087 6500 6111 6502
rect 6167 6500 6173 6502
rect 5865 6491 6173 6500
rect 5172 6452 5224 6458
rect 5172 6394 5224 6400
rect 5205 6012 5513 6021
rect 5205 6010 5211 6012
rect 5267 6010 5291 6012
rect 5347 6010 5371 6012
rect 5427 6010 5451 6012
rect 5507 6010 5513 6012
rect 5267 5958 5269 6010
rect 5449 5958 5451 6010
rect 5205 5956 5211 5958
rect 5267 5956 5291 5958
rect 5347 5956 5371 5958
rect 5427 5956 5451 5958
rect 5507 5956 5513 5958
rect 5205 5947 5513 5956
rect 5080 5908 5132 5914
rect 5000 5868 5080 5896
rect 4896 5024 4948 5030
rect 4896 4966 4948 4972
rect 4908 4826 4936 4966
rect 4896 4820 4948 4826
rect 4896 4762 4948 4768
rect 4804 4684 4856 4690
rect 4804 4626 4856 4632
rect 4580 4576 4752 4604
rect 4528 4558 4580 4564
rect 4160 4480 4212 4486
rect 4160 4422 4212 4428
rect 4436 4480 4488 4486
rect 4436 4422 4488 4428
rect 4163 4380 4471 4389
rect 4163 4378 4169 4380
rect 4225 4378 4249 4380
rect 4305 4378 4329 4380
rect 4385 4378 4409 4380
rect 4465 4378 4471 4380
rect 4225 4326 4227 4378
rect 4407 4326 4409 4378
rect 4163 4324 4169 4326
rect 4225 4324 4249 4326
rect 4305 4324 4329 4326
rect 4385 4324 4409 4326
rect 4465 4324 4471 4326
rect 4163 4315 4471 4324
rect 4436 4208 4488 4214
rect 4434 4176 4436 4185
rect 4488 4176 4490 4185
rect 4434 4111 4490 4120
rect 4160 4004 4212 4010
rect 4160 3946 4212 3952
rect 3896 3862 4108 3890
rect 3503 3836 3811 3845
rect 3503 3834 3509 3836
rect 3565 3834 3589 3836
rect 3645 3834 3669 3836
rect 3725 3834 3749 3836
rect 3805 3834 3811 3836
rect 3565 3782 3567 3834
rect 3747 3782 3749 3834
rect 3503 3780 3509 3782
rect 3565 3780 3589 3782
rect 3645 3780 3669 3782
rect 3725 3780 3749 3782
rect 3805 3780 3811 3782
rect 3503 3771 3811 3780
rect 3436 3590 3556 3618
rect 3528 3398 3556 3590
rect 4080 3534 4108 3862
rect 4172 3738 4200 3946
rect 4160 3732 4212 3738
rect 4160 3674 4212 3680
rect 4540 3534 4568 4558
rect 4712 4480 4764 4486
rect 4712 4422 4764 4428
rect 4620 4140 4672 4146
rect 4620 4082 4672 4088
rect 4068 3528 4120 3534
rect 4068 3470 4120 3476
rect 4528 3528 4580 3534
rect 4528 3470 4580 3476
rect 3516 3392 3568 3398
rect 3516 3334 3568 3340
rect 3528 3058 3556 3334
rect 4163 3292 4471 3301
rect 4163 3290 4169 3292
rect 4225 3290 4249 3292
rect 4305 3290 4329 3292
rect 4385 3290 4409 3292
rect 4465 3290 4471 3292
rect 4225 3238 4227 3290
rect 4407 3238 4409 3290
rect 4163 3236 4169 3238
rect 4225 3236 4249 3238
rect 4305 3236 4329 3238
rect 4385 3236 4409 3238
rect 4465 3236 4471 3238
rect 4163 3227 4471 3236
rect 3516 3052 3568 3058
rect 3516 2994 3568 3000
rect 4540 2990 4568 3470
rect 4528 2984 4580 2990
rect 4528 2926 4580 2932
rect 3503 2748 3811 2757
rect 3503 2746 3509 2748
rect 3565 2746 3589 2748
rect 3645 2746 3669 2748
rect 3725 2746 3749 2748
rect 3805 2746 3811 2748
rect 3565 2694 3567 2746
rect 3747 2694 3749 2746
rect 3503 2692 3509 2694
rect 3565 2692 3589 2694
rect 3645 2692 3669 2694
rect 3725 2692 3749 2694
rect 3805 2692 3811 2694
rect 3503 2683 3811 2692
rect 4632 2650 4660 4082
rect 4724 3738 4752 4422
rect 4712 3732 4764 3738
rect 4712 3674 4764 3680
rect 4724 2650 4752 3674
rect 4816 3602 4844 4626
rect 4908 4486 4936 4762
rect 4896 4480 4948 4486
rect 4896 4422 4948 4428
rect 4896 4004 4948 4010
rect 4896 3946 4948 3952
rect 4804 3596 4856 3602
rect 4804 3538 4856 3544
rect 4620 2644 4672 2650
rect 4620 2586 4672 2592
rect 4712 2644 4764 2650
rect 4712 2586 4764 2592
rect 4816 2446 4844 3538
rect 4908 3194 4936 3946
rect 4896 3188 4948 3194
rect 4896 3130 4948 3136
rect 5000 3126 5028 5868
rect 5080 5850 5132 5856
rect 5865 5468 6173 5477
rect 5865 5466 5871 5468
rect 5927 5466 5951 5468
rect 6007 5466 6031 5468
rect 6087 5466 6111 5468
rect 6167 5466 6173 5468
rect 5927 5414 5929 5466
rect 6109 5414 6111 5466
rect 5865 5412 5871 5414
rect 5927 5412 5951 5414
rect 6007 5412 6031 5414
rect 6087 5412 6111 5414
rect 6167 5412 6173 5414
rect 5865 5403 6173 5412
rect 6288 5166 6316 6666
rect 6380 6458 6408 7278
rect 6368 6452 6420 6458
rect 6368 6394 6420 6400
rect 6656 6390 6684 7278
rect 6644 6384 6696 6390
rect 6644 6326 6696 6332
rect 6276 5160 6328 5166
rect 6276 5102 6328 5108
rect 5540 5024 5592 5030
rect 5540 4966 5592 4972
rect 5205 4924 5513 4933
rect 5205 4922 5211 4924
rect 5267 4922 5291 4924
rect 5347 4922 5371 4924
rect 5427 4922 5451 4924
rect 5507 4922 5513 4924
rect 5267 4870 5269 4922
rect 5449 4870 5451 4922
rect 5205 4868 5211 4870
rect 5267 4868 5291 4870
rect 5347 4868 5371 4870
rect 5427 4868 5451 4870
rect 5507 4868 5513 4870
rect 5205 4859 5513 4868
rect 5080 4616 5132 4622
rect 5080 4558 5132 4564
rect 5092 3516 5120 4558
rect 5264 4480 5316 4486
rect 5264 4422 5316 4428
rect 5276 4146 5304 4422
rect 5552 4146 5580 4966
rect 6288 4554 6316 5102
rect 6552 5024 6604 5030
rect 6552 4966 6604 4972
rect 5632 4548 5684 4554
rect 5632 4490 5684 4496
rect 6276 4548 6328 4554
rect 6276 4490 6328 4496
rect 5644 4282 5672 4490
rect 5865 4380 6173 4389
rect 5865 4378 5871 4380
rect 5927 4378 5951 4380
rect 6007 4378 6031 4380
rect 6087 4378 6111 4380
rect 6167 4378 6173 4380
rect 5927 4326 5929 4378
rect 6109 4326 6111 4378
rect 5865 4324 5871 4326
rect 5927 4324 5951 4326
rect 6007 4324 6031 4326
rect 6087 4324 6111 4326
rect 6167 4324 6173 4326
rect 5865 4315 6173 4324
rect 5632 4276 5684 4282
rect 5632 4218 5684 4224
rect 5630 4176 5686 4185
rect 5264 4140 5316 4146
rect 5264 4082 5316 4088
rect 5356 4140 5408 4146
rect 5356 4082 5408 4088
rect 5540 4140 5592 4146
rect 5630 4111 5632 4120
rect 5540 4082 5592 4088
rect 5684 4111 5686 4120
rect 5632 4082 5684 4088
rect 5368 3924 5396 4082
rect 5724 3936 5776 3942
rect 5368 3896 5580 3924
rect 5205 3836 5513 3845
rect 5205 3834 5211 3836
rect 5267 3834 5291 3836
rect 5347 3834 5371 3836
rect 5427 3834 5451 3836
rect 5507 3834 5513 3836
rect 5267 3782 5269 3834
rect 5449 3782 5451 3834
rect 5205 3780 5211 3782
rect 5267 3780 5291 3782
rect 5347 3780 5371 3782
rect 5427 3780 5451 3782
rect 5507 3780 5513 3782
rect 5205 3771 5513 3780
rect 5356 3732 5408 3738
rect 5552 3720 5580 3896
rect 5724 3878 5776 3884
rect 5408 3692 5580 3720
rect 5356 3674 5408 3680
rect 5736 3602 5764 3878
rect 5724 3596 5776 3602
rect 5724 3538 5776 3544
rect 5264 3528 5316 3534
rect 5092 3488 5264 3516
rect 4988 3120 5040 3126
rect 4988 3062 5040 3068
rect 5092 2990 5120 3488
rect 5264 3470 5316 3476
rect 6288 3466 6316 4490
rect 6564 4078 6592 4966
rect 6656 4690 6684 6326
rect 6840 6304 6868 8026
rect 6920 7744 6972 7750
rect 6920 7686 6972 7692
rect 6932 7478 6960 7686
rect 6920 7472 6972 7478
rect 6920 7414 6972 7420
rect 6932 7342 6960 7414
rect 6920 7336 6972 7342
rect 6920 7278 6972 7284
rect 6907 7100 7215 7109
rect 6907 7098 6913 7100
rect 6969 7098 6993 7100
rect 7049 7098 7073 7100
rect 7129 7098 7153 7100
rect 7209 7098 7215 7100
rect 6969 7046 6971 7098
rect 7151 7046 7153 7098
rect 6907 7044 6913 7046
rect 6969 7044 6993 7046
rect 7049 7044 7073 7046
rect 7129 7044 7153 7046
rect 7209 7044 7215 7046
rect 6907 7035 7215 7044
rect 7300 6474 7328 8298
rect 7392 6662 7420 8434
rect 7472 8424 7524 8430
rect 7472 8366 7524 8372
rect 7484 7886 7512 8366
rect 7472 7880 7524 7886
rect 7472 7822 7524 7828
rect 7567 7644 7875 7653
rect 7567 7642 7573 7644
rect 7629 7642 7653 7644
rect 7709 7642 7733 7644
rect 7789 7642 7813 7644
rect 7869 7642 7875 7644
rect 7629 7590 7631 7642
rect 7811 7590 7813 7642
rect 7567 7588 7573 7590
rect 7629 7588 7653 7590
rect 7709 7588 7733 7590
rect 7789 7588 7813 7590
rect 7869 7588 7875 7590
rect 7567 7579 7875 7588
rect 7944 7546 7972 8758
rect 8022 8735 8078 8744
rect 8024 7744 8076 7750
rect 8022 7712 8024 7721
rect 8076 7712 8078 7721
rect 8022 7647 8078 7656
rect 7932 7540 7984 7546
rect 7932 7482 7984 7488
rect 7472 7404 7524 7410
rect 7472 7346 7524 7352
rect 7484 7002 7512 7346
rect 7472 6996 7524 7002
rect 7472 6938 7524 6944
rect 7380 6656 7432 6662
rect 7380 6598 7432 6604
rect 7116 6446 7328 6474
rect 7116 6390 7144 6446
rect 7104 6384 7156 6390
rect 7104 6326 7156 6332
rect 7484 6322 7512 6938
rect 8022 6624 8078 6633
rect 7567 6556 7875 6565
rect 8022 6559 8078 6568
rect 7567 6554 7573 6556
rect 7629 6554 7653 6556
rect 7709 6554 7733 6556
rect 7789 6554 7813 6556
rect 7869 6554 7875 6556
rect 7629 6502 7631 6554
rect 7811 6502 7813 6554
rect 7567 6500 7573 6502
rect 7629 6500 7653 6502
rect 7709 6500 7733 6502
rect 7789 6500 7813 6502
rect 7869 6500 7875 6502
rect 7567 6491 7875 6500
rect 8036 6458 8064 6559
rect 8024 6452 8076 6458
rect 8024 6394 8076 6400
rect 6920 6316 6972 6322
rect 6840 6276 6920 6304
rect 6920 6258 6972 6264
rect 7472 6316 7524 6322
rect 7472 6258 7524 6264
rect 6907 6012 7215 6021
rect 6907 6010 6913 6012
rect 6969 6010 6993 6012
rect 7049 6010 7073 6012
rect 7129 6010 7153 6012
rect 7209 6010 7215 6012
rect 6969 5958 6971 6010
rect 7151 5958 7153 6010
rect 6907 5956 6913 5958
rect 6969 5956 6993 5958
rect 7049 5956 7073 5958
rect 7129 5956 7153 5958
rect 7209 5956 7215 5958
rect 6907 5947 7215 5956
rect 8024 5568 8076 5574
rect 8022 5536 8024 5545
rect 8076 5536 8078 5545
rect 7567 5468 7875 5477
rect 8022 5471 8078 5480
rect 7567 5466 7573 5468
rect 7629 5466 7653 5468
rect 7709 5466 7733 5468
rect 7789 5466 7813 5468
rect 7869 5466 7875 5468
rect 7629 5414 7631 5466
rect 7811 5414 7813 5466
rect 7567 5412 7573 5414
rect 7629 5412 7653 5414
rect 7709 5412 7733 5414
rect 7789 5412 7813 5414
rect 7869 5412 7875 5414
rect 7567 5403 7875 5412
rect 7380 5228 7432 5234
rect 7380 5170 7432 5176
rect 6907 4924 7215 4933
rect 6907 4922 6913 4924
rect 6969 4922 6993 4924
rect 7049 4922 7073 4924
rect 7129 4922 7153 4924
rect 7209 4922 7215 4924
rect 6969 4870 6971 4922
rect 7151 4870 7153 4922
rect 6907 4868 6913 4870
rect 6969 4868 6993 4870
rect 7049 4868 7073 4870
rect 7129 4868 7153 4870
rect 7209 4868 7215 4870
rect 6907 4859 7215 4868
rect 6644 4684 6696 4690
rect 6644 4626 6696 4632
rect 6828 4684 6880 4690
rect 6828 4626 6880 4632
rect 6656 4078 6684 4626
rect 6840 4146 6868 4626
rect 7392 4486 7420 5170
rect 7380 4480 7432 4486
rect 8024 4480 8076 4486
rect 7380 4422 7432 4428
rect 8022 4448 8024 4457
rect 8076 4448 8078 4457
rect 6828 4140 6880 4146
rect 6828 4082 6880 4088
rect 6552 4072 6604 4078
rect 6552 4014 6604 4020
rect 6644 4072 6696 4078
rect 6644 4014 6696 4020
rect 5632 3460 5684 3466
rect 5632 3402 5684 3408
rect 6276 3460 6328 3466
rect 6276 3402 6328 3408
rect 5644 3194 5672 3402
rect 5865 3292 6173 3301
rect 5865 3290 5871 3292
rect 5927 3290 5951 3292
rect 6007 3290 6031 3292
rect 6087 3290 6111 3292
rect 6167 3290 6173 3292
rect 5927 3238 5929 3290
rect 6109 3238 6111 3290
rect 5865 3236 5871 3238
rect 5927 3236 5951 3238
rect 6007 3236 6031 3238
rect 6087 3236 6111 3238
rect 6167 3236 6173 3238
rect 5865 3227 6173 3236
rect 5632 3188 5684 3194
rect 5632 3130 5684 3136
rect 6564 2990 6592 4014
rect 6656 3058 6684 4014
rect 7288 3936 7340 3942
rect 7288 3878 7340 3884
rect 6907 3836 7215 3845
rect 6907 3834 6913 3836
rect 6969 3834 6993 3836
rect 7049 3834 7073 3836
rect 7129 3834 7153 3836
rect 7209 3834 7215 3836
rect 6969 3782 6971 3834
rect 7151 3782 7153 3834
rect 6907 3780 6913 3782
rect 6969 3780 6993 3782
rect 7049 3780 7073 3782
rect 7129 3780 7153 3782
rect 7209 3780 7215 3782
rect 6907 3771 7215 3780
rect 7300 3534 7328 3878
rect 7288 3528 7340 3534
rect 7288 3470 7340 3476
rect 6920 3392 6972 3398
rect 6920 3334 6972 3340
rect 6932 3194 6960 3334
rect 6920 3188 6972 3194
rect 6920 3130 6972 3136
rect 7392 3058 7420 4422
rect 7567 4380 7875 4389
rect 8022 4383 8078 4392
rect 7567 4378 7573 4380
rect 7629 4378 7653 4380
rect 7709 4378 7733 4380
rect 7789 4378 7813 4380
rect 7869 4378 7875 4380
rect 7629 4326 7631 4378
rect 7811 4326 7813 4378
rect 7567 4324 7573 4326
rect 7629 4324 7653 4326
rect 7709 4324 7733 4326
rect 7789 4324 7813 4326
rect 7869 4324 7875 4326
rect 7567 4315 7875 4324
rect 8024 3392 8076 3398
rect 8022 3360 8024 3369
rect 8076 3360 8078 3369
rect 7567 3292 7875 3301
rect 8022 3295 8078 3304
rect 7567 3290 7573 3292
rect 7629 3290 7653 3292
rect 7709 3290 7733 3292
rect 7789 3290 7813 3292
rect 7869 3290 7875 3292
rect 7629 3238 7631 3290
rect 7811 3238 7813 3290
rect 7567 3236 7573 3238
rect 7629 3236 7653 3238
rect 7709 3236 7733 3238
rect 7789 3236 7813 3238
rect 7869 3236 7875 3238
rect 7567 3227 7875 3236
rect 6644 3052 6696 3058
rect 6644 2994 6696 3000
rect 7380 3052 7432 3058
rect 7380 2994 7432 3000
rect 5080 2984 5132 2990
rect 5080 2926 5132 2932
rect 6552 2984 6604 2990
rect 6552 2926 6604 2932
rect 7288 2916 7340 2922
rect 7288 2858 7340 2864
rect 5205 2748 5513 2757
rect 5205 2746 5211 2748
rect 5267 2746 5291 2748
rect 5347 2746 5371 2748
rect 5427 2746 5451 2748
rect 5507 2746 5513 2748
rect 5267 2694 5269 2746
rect 5449 2694 5451 2746
rect 5205 2692 5211 2694
rect 5267 2692 5291 2694
rect 5347 2692 5371 2694
rect 5427 2692 5451 2694
rect 5507 2692 5513 2694
rect 5205 2683 5513 2692
rect 6907 2748 7215 2757
rect 6907 2746 6913 2748
rect 6969 2746 6993 2748
rect 7049 2746 7073 2748
rect 7129 2746 7153 2748
rect 7209 2746 7215 2748
rect 6969 2694 6971 2746
rect 7151 2694 7153 2746
rect 6907 2692 6913 2694
rect 6969 2692 6993 2694
rect 7049 2692 7073 2694
rect 7129 2692 7153 2694
rect 7209 2692 7215 2694
rect 6907 2683 7215 2692
rect 7300 2446 7328 2858
rect 8024 2848 8076 2854
rect 8024 2790 8076 2796
rect 3332 2440 3384 2446
rect 3332 2382 3384 2388
rect 4804 2440 4856 2446
rect 4804 2382 4856 2388
rect 7288 2440 7340 2446
rect 7288 2382 7340 2388
rect 6828 2304 6880 2310
rect 8036 2281 8064 2790
rect 6828 2246 6880 2252
rect 8022 2272 8078 2281
rect 4163 2204 4471 2213
rect 4163 2202 4169 2204
rect 4225 2202 4249 2204
rect 4305 2202 4329 2204
rect 4385 2202 4409 2204
rect 4465 2202 4471 2204
rect 4225 2150 4227 2202
rect 4407 2150 4409 2202
rect 4163 2148 4169 2150
rect 4225 2148 4249 2150
rect 4305 2148 4329 2150
rect 4385 2148 4409 2150
rect 4465 2148 4471 2150
rect 4163 2139 4471 2148
rect 5865 2204 6173 2213
rect 5865 2202 5871 2204
rect 5927 2202 5951 2204
rect 6007 2202 6031 2204
rect 6087 2202 6111 2204
rect 6167 2202 6173 2204
rect 5927 2150 5929 2202
rect 6109 2150 6111 2202
rect 5865 2148 5871 2150
rect 5927 2148 5951 2150
rect 6007 2148 6031 2150
rect 6087 2148 6111 2150
rect 6167 2148 6173 2150
rect 5865 2139 6173 2148
rect 1764 1694 2934 1718
rect 1764 1532 1804 1694
rect 2874 1532 2934 1694
rect 1764 1504 2934 1532
rect 6840 1193 6868 2246
rect 7567 2204 7875 2213
rect 8022 2207 8078 2216
rect 7567 2202 7573 2204
rect 7629 2202 7653 2204
rect 7709 2202 7733 2204
rect 7789 2202 7813 2204
rect 7869 2202 7875 2204
rect 7629 2150 7631 2202
rect 7811 2150 7813 2202
rect 7567 2148 7573 2150
rect 7629 2148 7653 2150
rect 7709 2148 7733 2150
rect 7789 2148 7813 2150
rect 7869 2148 7875 2150
rect 7567 2139 7875 2148
rect 6826 1184 6882 1193
rect 6826 1119 6882 1128
<< via2 >>
rect 6642 9832 6698 9888
rect 2467 8730 2523 8732
rect 2547 8730 2603 8732
rect 2627 8730 2683 8732
rect 2707 8730 2763 8732
rect 2467 8678 2513 8730
rect 2513 8678 2523 8730
rect 2547 8678 2577 8730
rect 2577 8678 2589 8730
rect 2589 8678 2603 8730
rect 2627 8678 2641 8730
rect 2641 8678 2653 8730
rect 2653 8678 2683 8730
rect 2707 8678 2717 8730
rect 2717 8678 2763 8730
rect 2467 8676 2523 8678
rect 2547 8676 2603 8678
rect 2627 8676 2683 8678
rect 2707 8676 2763 8678
rect 4169 8730 4225 8732
rect 4249 8730 4305 8732
rect 4329 8730 4385 8732
rect 4409 8730 4465 8732
rect 4169 8678 4215 8730
rect 4215 8678 4225 8730
rect 4249 8678 4279 8730
rect 4279 8678 4291 8730
rect 4291 8678 4305 8730
rect 4329 8678 4343 8730
rect 4343 8678 4355 8730
rect 4355 8678 4385 8730
rect 4409 8678 4419 8730
rect 4419 8678 4465 8730
rect 4169 8676 4225 8678
rect 4249 8676 4305 8678
rect 4329 8676 4385 8678
rect 4409 8676 4465 8678
rect 5871 8730 5927 8732
rect 5951 8730 6007 8732
rect 6031 8730 6087 8732
rect 6111 8730 6167 8732
rect 5871 8678 5917 8730
rect 5917 8678 5927 8730
rect 5951 8678 5981 8730
rect 5981 8678 5993 8730
rect 5993 8678 6007 8730
rect 6031 8678 6045 8730
rect 6045 8678 6057 8730
rect 6057 8678 6087 8730
rect 6111 8678 6121 8730
rect 6121 8678 6167 8730
rect 5871 8676 5927 8678
rect 5951 8676 6007 8678
rect 6031 8676 6087 8678
rect 6111 8676 6167 8678
rect 7573 8730 7629 8732
rect 7653 8730 7709 8732
rect 7733 8730 7789 8732
rect 7813 8730 7869 8732
rect 7573 8678 7619 8730
rect 7619 8678 7629 8730
rect 7653 8678 7683 8730
rect 7683 8678 7695 8730
rect 7695 8678 7709 8730
rect 7733 8678 7747 8730
rect 7747 8678 7759 8730
rect 7759 8678 7789 8730
rect 7813 8678 7823 8730
rect 7823 8678 7869 8730
rect 7573 8676 7629 8678
rect 7653 8676 7709 8678
rect 7733 8676 7789 8678
rect 7813 8676 7869 8678
rect 1807 8186 1863 8188
rect 1887 8186 1943 8188
rect 1967 8186 2023 8188
rect 2047 8186 2103 8188
rect 1807 8134 1853 8186
rect 1853 8134 1863 8186
rect 1887 8134 1917 8186
rect 1917 8134 1929 8186
rect 1929 8134 1943 8186
rect 1967 8134 1981 8186
rect 1981 8134 1993 8186
rect 1993 8134 2023 8186
rect 2047 8134 2057 8186
rect 2057 8134 2103 8186
rect 1807 8132 1863 8134
rect 1887 8132 1943 8134
rect 1967 8132 2023 8134
rect 2047 8132 2103 8134
rect 1807 7098 1863 7100
rect 1887 7098 1943 7100
rect 1967 7098 2023 7100
rect 2047 7098 2103 7100
rect 1807 7046 1853 7098
rect 1853 7046 1863 7098
rect 1887 7046 1917 7098
rect 1917 7046 1929 7098
rect 1929 7046 1943 7098
rect 1967 7046 1981 7098
rect 1981 7046 1993 7098
rect 1993 7046 2023 7098
rect 2047 7046 2057 7098
rect 2057 7046 2103 7098
rect 1807 7044 1863 7046
rect 1887 7044 1943 7046
rect 1967 7044 2023 7046
rect 2047 7044 2103 7046
rect 3509 8186 3565 8188
rect 3589 8186 3645 8188
rect 3669 8186 3725 8188
rect 3749 8186 3805 8188
rect 3509 8134 3555 8186
rect 3555 8134 3565 8186
rect 3589 8134 3619 8186
rect 3619 8134 3631 8186
rect 3631 8134 3645 8186
rect 3669 8134 3683 8186
rect 3683 8134 3695 8186
rect 3695 8134 3725 8186
rect 3749 8134 3759 8186
rect 3759 8134 3805 8186
rect 3509 8132 3565 8134
rect 3589 8132 3645 8134
rect 3669 8132 3725 8134
rect 3749 8132 3805 8134
rect 2467 7642 2523 7644
rect 2547 7642 2603 7644
rect 2627 7642 2683 7644
rect 2707 7642 2763 7644
rect 2467 7590 2513 7642
rect 2513 7590 2523 7642
rect 2547 7590 2577 7642
rect 2577 7590 2589 7642
rect 2589 7590 2603 7642
rect 2627 7590 2641 7642
rect 2641 7590 2653 7642
rect 2653 7590 2683 7642
rect 2707 7590 2717 7642
rect 2717 7590 2763 7642
rect 2467 7588 2523 7590
rect 2547 7588 2603 7590
rect 2627 7588 2683 7590
rect 2707 7588 2763 7590
rect 2467 6554 2523 6556
rect 2547 6554 2603 6556
rect 2627 6554 2683 6556
rect 2707 6554 2763 6556
rect 2467 6502 2513 6554
rect 2513 6502 2523 6554
rect 2547 6502 2577 6554
rect 2577 6502 2589 6554
rect 2589 6502 2603 6554
rect 2627 6502 2641 6554
rect 2641 6502 2653 6554
rect 2653 6502 2683 6554
rect 2707 6502 2717 6554
rect 2717 6502 2763 6554
rect 2467 6500 2523 6502
rect 2547 6500 2603 6502
rect 2627 6500 2683 6502
rect 2707 6500 2763 6502
rect 1807 6010 1863 6012
rect 1887 6010 1943 6012
rect 1967 6010 2023 6012
rect 2047 6010 2103 6012
rect 1807 5958 1853 6010
rect 1853 5958 1863 6010
rect 1887 5958 1917 6010
rect 1917 5958 1929 6010
rect 1929 5958 1943 6010
rect 1967 5958 1981 6010
rect 1981 5958 1993 6010
rect 1993 5958 2023 6010
rect 2047 5958 2057 6010
rect 2057 5958 2103 6010
rect 1807 5956 1863 5958
rect 1887 5956 1943 5958
rect 1967 5956 2023 5958
rect 2047 5956 2103 5958
rect 4169 7642 4225 7644
rect 4249 7642 4305 7644
rect 4329 7642 4385 7644
rect 4409 7642 4465 7644
rect 4169 7590 4215 7642
rect 4215 7590 4225 7642
rect 4249 7590 4279 7642
rect 4279 7590 4291 7642
rect 4291 7590 4305 7642
rect 4329 7590 4343 7642
rect 4343 7590 4355 7642
rect 4355 7590 4385 7642
rect 4409 7590 4419 7642
rect 4419 7590 4465 7642
rect 4169 7588 4225 7590
rect 4249 7588 4305 7590
rect 4329 7588 4385 7590
rect 4409 7588 4465 7590
rect 4434 7404 4490 7440
rect 4434 7384 4436 7404
rect 4436 7384 4488 7404
rect 4488 7384 4490 7404
rect 2467 5466 2523 5468
rect 2547 5466 2603 5468
rect 2627 5466 2683 5468
rect 2707 5466 2763 5468
rect 2467 5414 2513 5466
rect 2513 5414 2523 5466
rect 2547 5414 2577 5466
rect 2577 5414 2589 5466
rect 2589 5414 2603 5466
rect 2627 5414 2641 5466
rect 2641 5414 2653 5466
rect 2653 5414 2683 5466
rect 2707 5414 2717 5466
rect 2717 5414 2763 5466
rect 2467 5412 2523 5414
rect 2547 5412 2603 5414
rect 2627 5412 2683 5414
rect 2707 5412 2763 5414
rect 1807 4922 1863 4924
rect 1887 4922 1943 4924
rect 1967 4922 2023 4924
rect 2047 4922 2103 4924
rect 1807 4870 1853 4922
rect 1853 4870 1863 4922
rect 1887 4870 1917 4922
rect 1917 4870 1929 4922
rect 1929 4870 1943 4922
rect 1967 4870 1981 4922
rect 1981 4870 1993 4922
rect 1993 4870 2023 4922
rect 2047 4870 2057 4922
rect 2057 4870 2103 4922
rect 1807 4868 1863 4870
rect 1887 4868 1943 4870
rect 1967 4868 2023 4870
rect 2047 4868 2103 4870
rect 2467 4378 2523 4380
rect 2547 4378 2603 4380
rect 2627 4378 2683 4380
rect 2707 4378 2763 4380
rect 2467 4326 2513 4378
rect 2513 4326 2523 4378
rect 2547 4326 2577 4378
rect 2577 4326 2589 4378
rect 2589 4326 2603 4378
rect 2627 4326 2641 4378
rect 2641 4326 2653 4378
rect 2653 4326 2683 4378
rect 2707 4326 2717 4378
rect 2717 4326 2763 4378
rect 2467 4324 2523 4326
rect 2547 4324 2603 4326
rect 2627 4324 2683 4326
rect 2707 4324 2763 4326
rect 1807 3834 1863 3836
rect 1887 3834 1943 3836
rect 1967 3834 2023 3836
rect 2047 3834 2103 3836
rect 1807 3782 1853 3834
rect 1853 3782 1863 3834
rect 1887 3782 1917 3834
rect 1917 3782 1929 3834
rect 1929 3782 1943 3834
rect 1967 3782 1981 3834
rect 1981 3782 1993 3834
rect 1993 3782 2023 3834
rect 2047 3782 2057 3834
rect 2057 3782 2103 3834
rect 1807 3780 1863 3782
rect 1887 3780 1943 3782
rect 1967 3780 2023 3782
rect 2047 3780 2103 3782
rect 2467 3290 2523 3292
rect 2547 3290 2603 3292
rect 2627 3290 2683 3292
rect 2707 3290 2763 3292
rect 2467 3238 2513 3290
rect 2513 3238 2523 3290
rect 2547 3238 2577 3290
rect 2577 3238 2589 3290
rect 2589 3238 2603 3290
rect 2627 3238 2641 3290
rect 2641 3238 2653 3290
rect 2653 3238 2683 3290
rect 2707 3238 2717 3290
rect 2717 3238 2763 3290
rect 2467 3236 2523 3238
rect 2547 3236 2603 3238
rect 2627 3236 2683 3238
rect 2707 3236 2763 3238
rect 1807 2746 1863 2748
rect 1887 2746 1943 2748
rect 1967 2746 2023 2748
rect 2047 2746 2103 2748
rect 1807 2694 1853 2746
rect 1853 2694 1863 2746
rect 1887 2694 1917 2746
rect 1917 2694 1929 2746
rect 1929 2694 1943 2746
rect 1967 2694 1981 2746
rect 1981 2694 1993 2746
rect 1993 2694 2023 2746
rect 2047 2694 2057 2746
rect 2057 2694 2103 2746
rect 1807 2692 1863 2694
rect 1887 2692 1943 2694
rect 1967 2692 2023 2694
rect 2047 2692 2103 2694
rect 2467 2202 2523 2204
rect 2547 2202 2603 2204
rect 2627 2202 2683 2204
rect 2707 2202 2763 2204
rect 2467 2150 2513 2202
rect 2513 2150 2523 2202
rect 2547 2150 2577 2202
rect 2577 2150 2589 2202
rect 2589 2150 2603 2202
rect 2627 2150 2641 2202
rect 2641 2150 2653 2202
rect 2653 2150 2683 2202
rect 2707 2150 2717 2202
rect 2717 2150 2763 2202
rect 2467 2148 2523 2150
rect 2547 2148 2603 2150
rect 2627 2148 2683 2150
rect 2707 2148 2763 2150
rect 3509 7098 3565 7100
rect 3589 7098 3645 7100
rect 3669 7098 3725 7100
rect 3749 7098 3805 7100
rect 3509 7046 3555 7098
rect 3555 7046 3565 7098
rect 3589 7046 3619 7098
rect 3619 7046 3631 7098
rect 3631 7046 3645 7098
rect 3669 7046 3683 7098
rect 3683 7046 3695 7098
rect 3695 7046 3725 7098
rect 3749 7046 3759 7098
rect 3759 7046 3805 7098
rect 3509 7044 3565 7046
rect 3589 7044 3645 7046
rect 3669 7044 3725 7046
rect 3749 7044 3805 7046
rect 4169 6554 4225 6556
rect 4249 6554 4305 6556
rect 4329 6554 4385 6556
rect 4409 6554 4465 6556
rect 4169 6502 4215 6554
rect 4215 6502 4225 6554
rect 4249 6502 4279 6554
rect 4279 6502 4291 6554
rect 4291 6502 4305 6554
rect 4329 6502 4343 6554
rect 4343 6502 4355 6554
rect 4355 6502 4385 6554
rect 4409 6502 4419 6554
rect 4419 6502 4465 6554
rect 4169 6500 4225 6502
rect 4249 6500 4305 6502
rect 4329 6500 4385 6502
rect 4409 6500 4465 6502
rect 3509 6010 3565 6012
rect 3589 6010 3645 6012
rect 3669 6010 3725 6012
rect 3749 6010 3805 6012
rect 3509 5958 3555 6010
rect 3555 5958 3565 6010
rect 3589 5958 3619 6010
rect 3619 5958 3631 6010
rect 3631 5958 3645 6010
rect 3669 5958 3683 6010
rect 3683 5958 3695 6010
rect 3695 5958 3725 6010
rect 3749 5958 3759 6010
rect 3759 5958 3805 6010
rect 3509 5956 3565 5958
rect 3589 5956 3645 5958
rect 3669 5956 3725 5958
rect 3749 5956 3805 5958
rect 4169 5466 4225 5468
rect 4249 5466 4305 5468
rect 4329 5466 4385 5468
rect 4409 5466 4465 5468
rect 4169 5414 4215 5466
rect 4215 5414 4225 5466
rect 4249 5414 4279 5466
rect 4279 5414 4291 5466
rect 4291 5414 4305 5466
rect 4329 5414 4343 5466
rect 4343 5414 4355 5466
rect 4355 5414 4385 5466
rect 4409 5414 4419 5466
rect 4419 5414 4465 5466
rect 4169 5412 4225 5414
rect 4249 5412 4305 5414
rect 4329 5412 4385 5414
rect 4409 5412 4465 5414
rect 3509 4922 3565 4924
rect 3589 4922 3645 4924
rect 3669 4922 3725 4924
rect 3749 4922 3805 4924
rect 3509 4870 3555 4922
rect 3555 4870 3565 4922
rect 3589 4870 3619 4922
rect 3619 4870 3631 4922
rect 3631 4870 3645 4922
rect 3669 4870 3683 4922
rect 3683 4870 3695 4922
rect 3695 4870 3725 4922
rect 3749 4870 3759 4922
rect 3759 4870 3805 4922
rect 3509 4868 3565 4870
rect 3589 4868 3645 4870
rect 3669 4868 3725 4870
rect 3749 4868 3805 4870
rect 5211 8186 5267 8188
rect 5291 8186 5347 8188
rect 5371 8186 5427 8188
rect 5451 8186 5507 8188
rect 5211 8134 5257 8186
rect 5257 8134 5267 8186
rect 5291 8134 5321 8186
rect 5321 8134 5333 8186
rect 5333 8134 5347 8186
rect 5371 8134 5385 8186
rect 5385 8134 5397 8186
rect 5397 8134 5427 8186
rect 5451 8134 5461 8186
rect 5461 8134 5507 8186
rect 5211 8132 5267 8134
rect 5291 8132 5347 8134
rect 5371 8132 5427 8134
rect 5451 8132 5507 8134
rect 6913 8186 6969 8188
rect 6993 8186 7049 8188
rect 7073 8186 7129 8188
rect 7153 8186 7209 8188
rect 6913 8134 6959 8186
rect 6959 8134 6969 8186
rect 6993 8134 7023 8186
rect 7023 8134 7035 8186
rect 7035 8134 7049 8186
rect 7073 8134 7087 8186
rect 7087 8134 7099 8186
rect 7099 8134 7129 8186
rect 7153 8134 7163 8186
rect 7163 8134 7209 8186
rect 6913 8132 6969 8134
rect 6993 8132 7049 8134
rect 7073 8132 7129 8134
rect 7153 8132 7209 8134
rect 5262 7384 5318 7440
rect 5211 7098 5267 7100
rect 5291 7098 5347 7100
rect 5371 7098 5427 7100
rect 5451 7098 5507 7100
rect 5211 7046 5257 7098
rect 5257 7046 5267 7098
rect 5291 7046 5321 7098
rect 5321 7046 5333 7098
rect 5333 7046 5347 7098
rect 5371 7046 5385 7098
rect 5385 7046 5397 7098
rect 5397 7046 5427 7098
rect 5451 7046 5461 7098
rect 5461 7046 5507 7098
rect 5211 7044 5267 7046
rect 5291 7044 5347 7046
rect 5371 7044 5427 7046
rect 5451 7044 5507 7046
rect 5871 7642 5927 7644
rect 5951 7642 6007 7644
rect 6031 7642 6087 7644
rect 6111 7642 6167 7644
rect 5871 7590 5917 7642
rect 5917 7590 5927 7642
rect 5951 7590 5981 7642
rect 5981 7590 5993 7642
rect 5993 7590 6007 7642
rect 6031 7590 6045 7642
rect 6045 7590 6057 7642
rect 6057 7590 6087 7642
rect 6111 7590 6121 7642
rect 6121 7590 6167 7642
rect 5871 7588 5927 7590
rect 5951 7588 6007 7590
rect 6031 7588 6087 7590
rect 6111 7588 6167 7590
rect 5871 6554 5927 6556
rect 5951 6554 6007 6556
rect 6031 6554 6087 6556
rect 6111 6554 6167 6556
rect 5871 6502 5917 6554
rect 5917 6502 5927 6554
rect 5951 6502 5981 6554
rect 5981 6502 5993 6554
rect 5993 6502 6007 6554
rect 6031 6502 6045 6554
rect 6045 6502 6057 6554
rect 6057 6502 6087 6554
rect 6111 6502 6121 6554
rect 6121 6502 6167 6554
rect 5871 6500 5927 6502
rect 5951 6500 6007 6502
rect 6031 6500 6087 6502
rect 6111 6500 6167 6502
rect 5211 6010 5267 6012
rect 5291 6010 5347 6012
rect 5371 6010 5427 6012
rect 5451 6010 5507 6012
rect 5211 5958 5257 6010
rect 5257 5958 5267 6010
rect 5291 5958 5321 6010
rect 5321 5958 5333 6010
rect 5333 5958 5347 6010
rect 5371 5958 5385 6010
rect 5385 5958 5397 6010
rect 5397 5958 5427 6010
rect 5451 5958 5461 6010
rect 5461 5958 5507 6010
rect 5211 5956 5267 5958
rect 5291 5956 5347 5958
rect 5371 5956 5427 5958
rect 5451 5956 5507 5958
rect 4169 4378 4225 4380
rect 4249 4378 4305 4380
rect 4329 4378 4385 4380
rect 4409 4378 4465 4380
rect 4169 4326 4215 4378
rect 4215 4326 4225 4378
rect 4249 4326 4279 4378
rect 4279 4326 4291 4378
rect 4291 4326 4305 4378
rect 4329 4326 4343 4378
rect 4343 4326 4355 4378
rect 4355 4326 4385 4378
rect 4409 4326 4419 4378
rect 4419 4326 4465 4378
rect 4169 4324 4225 4326
rect 4249 4324 4305 4326
rect 4329 4324 4385 4326
rect 4409 4324 4465 4326
rect 4434 4156 4436 4176
rect 4436 4156 4488 4176
rect 4488 4156 4490 4176
rect 4434 4120 4490 4156
rect 3509 3834 3565 3836
rect 3589 3834 3645 3836
rect 3669 3834 3725 3836
rect 3749 3834 3805 3836
rect 3509 3782 3555 3834
rect 3555 3782 3565 3834
rect 3589 3782 3619 3834
rect 3619 3782 3631 3834
rect 3631 3782 3645 3834
rect 3669 3782 3683 3834
rect 3683 3782 3695 3834
rect 3695 3782 3725 3834
rect 3749 3782 3759 3834
rect 3759 3782 3805 3834
rect 3509 3780 3565 3782
rect 3589 3780 3645 3782
rect 3669 3780 3725 3782
rect 3749 3780 3805 3782
rect 4169 3290 4225 3292
rect 4249 3290 4305 3292
rect 4329 3290 4385 3292
rect 4409 3290 4465 3292
rect 4169 3238 4215 3290
rect 4215 3238 4225 3290
rect 4249 3238 4279 3290
rect 4279 3238 4291 3290
rect 4291 3238 4305 3290
rect 4329 3238 4343 3290
rect 4343 3238 4355 3290
rect 4355 3238 4385 3290
rect 4409 3238 4419 3290
rect 4419 3238 4465 3290
rect 4169 3236 4225 3238
rect 4249 3236 4305 3238
rect 4329 3236 4385 3238
rect 4409 3236 4465 3238
rect 3509 2746 3565 2748
rect 3589 2746 3645 2748
rect 3669 2746 3725 2748
rect 3749 2746 3805 2748
rect 3509 2694 3555 2746
rect 3555 2694 3565 2746
rect 3589 2694 3619 2746
rect 3619 2694 3631 2746
rect 3631 2694 3645 2746
rect 3669 2694 3683 2746
rect 3683 2694 3695 2746
rect 3695 2694 3725 2746
rect 3749 2694 3759 2746
rect 3759 2694 3805 2746
rect 3509 2692 3565 2694
rect 3589 2692 3645 2694
rect 3669 2692 3725 2694
rect 3749 2692 3805 2694
rect 5871 5466 5927 5468
rect 5951 5466 6007 5468
rect 6031 5466 6087 5468
rect 6111 5466 6167 5468
rect 5871 5414 5917 5466
rect 5917 5414 5927 5466
rect 5951 5414 5981 5466
rect 5981 5414 5993 5466
rect 5993 5414 6007 5466
rect 6031 5414 6045 5466
rect 6045 5414 6057 5466
rect 6057 5414 6087 5466
rect 6111 5414 6121 5466
rect 6121 5414 6167 5466
rect 5871 5412 5927 5414
rect 5951 5412 6007 5414
rect 6031 5412 6087 5414
rect 6111 5412 6167 5414
rect 5211 4922 5267 4924
rect 5291 4922 5347 4924
rect 5371 4922 5427 4924
rect 5451 4922 5507 4924
rect 5211 4870 5257 4922
rect 5257 4870 5267 4922
rect 5291 4870 5321 4922
rect 5321 4870 5333 4922
rect 5333 4870 5347 4922
rect 5371 4870 5385 4922
rect 5385 4870 5397 4922
rect 5397 4870 5427 4922
rect 5451 4870 5461 4922
rect 5461 4870 5507 4922
rect 5211 4868 5267 4870
rect 5291 4868 5347 4870
rect 5371 4868 5427 4870
rect 5451 4868 5507 4870
rect 5871 4378 5927 4380
rect 5951 4378 6007 4380
rect 6031 4378 6087 4380
rect 6111 4378 6167 4380
rect 5871 4326 5917 4378
rect 5917 4326 5927 4378
rect 5951 4326 5981 4378
rect 5981 4326 5993 4378
rect 5993 4326 6007 4378
rect 6031 4326 6045 4378
rect 6045 4326 6057 4378
rect 6057 4326 6087 4378
rect 6111 4326 6121 4378
rect 6121 4326 6167 4378
rect 5871 4324 5927 4326
rect 5951 4324 6007 4326
rect 6031 4324 6087 4326
rect 6111 4324 6167 4326
rect 5630 4140 5686 4176
rect 5630 4120 5632 4140
rect 5632 4120 5684 4140
rect 5684 4120 5686 4140
rect 5211 3834 5267 3836
rect 5291 3834 5347 3836
rect 5371 3834 5427 3836
rect 5451 3834 5507 3836
rect 5211 3782 5257 3834
rect 5257 3782 5267 3834
rect 5291 3782 5321 3834
rect 5321 3782 5333 3834
rect 5333 3782 5347 3834
rect 5371 3782 5385 3834
rect 5385 3782 5397 3834
rect 5397 3782 5427 3834
rect 5451 3782 5461 3834
rect 5461 3782 5507 3834
rect 5211 3780 5267 3782
rect 5291 3780 5347 3782
rect 5371 3780 5427 3782
rect 5451 3780 5507 3782
rect 6913 7098 6969 7100
rect 6993 7098 7049 7100
rect 7073 7098 7129 7100
rect 7153 7098 7209 7100
rect 6913 7046 6959 7098
rect 6959 7046 6969 7098
rect 6993 7046 7023 7098
rect 7023 7046 7035 7098
rect 7035 7046 7049 7098
rect 7073 7046 7087 7098
rect 7087 7046 7099 7098
rect 7099 7046 7129 7098
rect 7153 7046 7163 7098
rect 7163 7046 7209 7098
rect 6913 7044 6969 7046
rect 6993 7044 7049 7046
rect 7073 7044 7129 7046
rect 7153 7044 7209 7046
rect 7573 7642 7629 7644
rect 7653 7642 7709 7644
rect 7733 7642 7789 7644
rect 7813 7642 7869 7644
rect 7573 7590 7619 7642
rect 7619 7590 7629 7642
rect 7653 7590 7683 7642
rect 7683 7590 7695 7642
rect 7695 7590 7709 7642
rect 7733 7590 7747 7642
rect 7747 7590 7759 7642
rect 7759 7590 7789 7642
rect 7813 7590 7823 7642
rect 7823 7590 7869 7642
rect 7573 7588 7629 7590
rect 7653 7588 7709 7590
rect 7733 7588 7789 7590
rect 7813 7588 7869 7590
rect 8022 8744 8078 8800
rect 8022 7692 8024 7712
rect 8024 7692 8076 7712
rect 8076 7692 8078 7712
rect 8022 7656 8078 7692
rect 8022 6568 8078 6624
rect 7573 6554 7629 6556
rect 7653 6554 7709 6556
rect 7733 6554 7789 6556
rect 7813 6554 7869 6556
rect 7573 6502 7619 6554
rect 7619 6502 7629 6554
rect 7653 6502 7683 6554
rect 7683 6502 7695 6554
rect 7695 6502 7709 6554
rect 7733 6502 7747 6554
rect 7747 6502 7759 6554
rect 7759 6502 7789 6554
rect 7813 6502 7823 6554
rect 7823 6502 7869 6554
rect 7573 6500 7629 6502
rect 7653 6500 7709 6502
rect 7733 6500 7789 6502
rect 7813 6500 7869 6502
rect 6913 6010 6969 6012
rect 6993 6010 7049 6012
rect 7073 6010 7129 6012
rect 7153 6010 7209 6012
rect 6913 5958 6959 6010
rect 6959 5958 6969 6010
rect 6993 5958 7023 6010
rect 7023 5958 7035 6010
rect 7035 5958 7049 6010
rect 7073 5958 7087 6010
rect 7087 5958 7099 6010
rect 7099 5958 7129 6010
rect 7153 5958 7163 6010
rect 7163 5958 7209 6010
rect 6913 5956 6969 5958
rect 6993 5956 7049 5958
rect 7073 5956 7129 5958
rect 7153 5956 7209 5958
rect 8022 5516 8024 5536
rect 8024 5516 8076 5536
rect 8076 5516 8078 5536
rect 8022 5480 8078 5516
rect 7573 5466 7629 5468
rect 7653 5466 7709 5468
rect 7733 5466 7789 5468
rect 7813 5466 7869 5468
rect 7573 5414 7619 5466
rect 7619 5414 7629 5466
rect 7653 5414 7683 5466
rect 7683 5414 7695 5466
rect 7695 5414 7709 5466
rect 7733 5414 7747 5466
rect 7747 5414 7759 5466
rect 7759 5414 7789 5466
rect 7813 5414 7823 5466
rect 7823 5414 7869 5466
rect 7573 5412 7629 5414
rect 7653 5412 7709 5414
rect 7733 5412 7789 5414
rect 7813 5412 7869 5414
rect 6913 4922 6969 4924
rect 6993 4922 7049 4924
rect 7073 4922 7129 4924
rect 7153 4922 7209 4924
rect 6913 4870 6959 4922
rect 6959 4870 6969 4922
rect 6993 4870 7023 4922
rect 7023 4870 7035 4922
rect 7035 4870 7049 4922
rect 7073 4870 7087 4922
rect 7087 4870 7099 4922
rect 7099 4870 7129 4922
rect 7153 4870 7163 4922
rect 7163 4870 7209 4922
rect 6913 4868 6969 4870
rect 6993 4868 7049 4870
rect 7073 4868 7129 4870
rect 7153 4868 7209 4870
rect 8022 4428 8024 4448
rect 8024 4428 8076 4448
rect 8076 4428 8078 4448
rect 5871 3290 5927 3292
rect 5951 3290 6007 3292
rect 6031 3290 6087 3292
rect 6111 3290 6167 3292
rect 5871 3238 5917 3290
rect 5917 3238 5927 3290
rect 5951 3238 5981 3290
rect 5981 3238 5993 3290
rect 5993 3238 6007 3290
rect 6031 3238 6045 3290
rect 6045 3238 6057 3290
rect 6057 3238 6087 3290
rect 6111 3238 6121 3290
rect 6121 3238 6167 3290
rect 5871 3236 5927 3238
rect 5951 3236 6007 3238
rect 6031 3236 6087 3238
rect 6111 3236 6167 3238
rect 6913 3834 6969 3836
rect 6993 3834 7049 3836
rect 7073 3834 7129 3836
rect 7153 3834 7209 3836
rect 6913 3782 6959 3834
rect 6959 3782 6969 3834
rect 6993 3782 7023 3834
rect 7023 3782 7035 3834
rect 7035 3782 7049 3834
rect 7073 3782 7087 3834
rect 7087 3782 7099 3834
rect 7099 3782 7129 3834
rect 7153 3782 7163 3834
rect 7163 3782 7209 3834
rect 6913 3780 6969 3782
rect 6993 3780 7049 3782
rect 7073 3780 7129 3782
rect 7153 3780 7209 3782
rect 8022 4392 8078 4428
rect 7573 4378 7629 4380
rect 7653 4378 7709 4380
rect 7733 4378 7789 4380
rect 7813 4378 7869 4380
rect 7573 4326 7619 4378
rect 7619 4326 7629 4378
rect 7653 4326 7683 4378
rect 7683 4326 7695 4378
rect 7695 4326 7709 4378
rect 7733 4326 7747 4378
rect 7747 4326 7759 4378
rect 7759 4326 7789 4378
rect 7813 4326 7823 4378
rect 7823 4326 7869 4378
rect 7573 4324 7629 4326
rect 7653 4324 7709 4326
rect 7733 4324 7789 4326
rect 7813 4324 7869 4326
rect 8022 3340 8024 3360
rect 8024 3340 8076 3360
rect 8076 3340 8078 3360
rect 8022 3304 8078 3340
rect 7573 3290 7629 3292
rect 7653 3290 7709 3292
rect 7733 3290 7789 3292
rect 7813 3290 7869 3292
rect 7573 3238 7619 3290
rect 7619 3238 7629 3290
rect 7653 3238 7683 3290
rect 7683 3238 7695 3290
rect 7695 3238 7709 3290
rect 7733 3238 7747 3290
rect 7747 3238 7759 3290
rect 7759 3238 7789 3290
rect 7813 3238 7823 3290
rect 7823 3238 7869 3290
rect 7573 3236 7629 3238
rect 7653 3236 7709 3238
rect 7733 3236 7789 3238
rect 7813 3236 7869 3238
rect 5211 2746 5267 2748
rect 5291 2746 5347 2748
rect 5371 2746 5427 2748
rect 5451 2746 5507 2748
rect 5211 2694 5257 2746
rect 5257 2694 5267 2746
rect 5291 2694 5321 2746
rect 5321 2694 5333 2746
rect 5333 2694 5347 2746
rect 5371 2694 5385 2746
rect 5385 2694 5397 2746
rect 5397 2694 5427 2746
rect 5451 2694 5461 2746
rect 5461 2694 5507 2746
rect 5211 2692 5267 2694
rect 5291 2692 5347 2694
rect 5371 2692 5427 2694
rect 5451 2692 5507 2694
rect 6913 2746 6969 2748
rect 6993 2746 7049 2748
rect 7073 2746 7129 2748
rect 7153 2746 7209 2748
rect 6913 2694 6959 2746
rect 6959 2694 6969 2746
rect 6993 2694 7023 2746
rect 7023 2694 7035 2746
rect 7035 2694 7049 2746
rect 7073 2694 7087 2746
rect 7087 2694 7099 2746
rect 7099 2694 7129 2746
rect 7153 2694 7163 2746
rect 7163 2694 7209 2746
rect 6913 2692 6969 2694
rect 6993 2692 7049 2694
rect 7073 2692 7129 2694
rect 7153 2692 7209 2694
rect 4169 2202 4225 2204
rect 4249 2202 4305 2204
rect 4329 2202 4385 2204
rect 4409 2202 4465 2204
rect 4169 2150 4215 2202
rect 4215 2150 4225 2202
rect 4249 2150 4279 2202
rect 4279 2150 4291 2202
rect 4291 2150 4305 2202
rect 4329 2150 4343 2202
rect 4343 2150 4355 2202
rect 4355 2150 4385 2202
rect 4409 2150 4419 2202
rect 4419 2150 4465 2202
rect 4169 2148 4225 2150
rect 4249 2148 4305 2150
rect 4329 2148 4385 2150
rect 4409 2148 4465 2150
rect 5871 2202 5927 2204
rect 5951 2202 6007 2204
rect 6031 2202 6087 2204
rect 6111 2202 6167 2204
rect 5871 2150 5917 2202
rect 5917 2150 5927 2202
rect 5951 2150 5981 2202
rect 5981 2150 5993 2202
rect 5993 2150 6007 2202
rect 6031 2150 6045 2202
rect 6045 2150 6057 2202
rect 6057 2150 6087 2202
rect 6111 2150 6121 2202
rect 6121 2150 6167 2202
rect 5871 2148 5927 2150
rect 5951 2148 6007 2150
rect 6031 2148 6087 2150
rect 6111 2148 6167 2150
rect 8022 2216 8078 2272
rect 7573 2202 7629 2204
rect 7653 2202 7709 2204
rect 7733 2202 7789 2204
rect 7813 2202 7869 2204
rect 7573 2150 7619 2202
rect 7619 2150 7629 2202
rect 7653 2150 7683 2202
rect 7683 2150 7695 2202
rect 7695 2150 7709 2202
rect 7733 2150 7747 2202
rect 7747 2150 7759 2202
rect 7759 2150 7789 2202
rect 7813 2150 7823 2202
rect 7823 2150 7869 2202
rect 7573 2148 7629 2150
rect 7653 2148 7709 2150
rect 7733 2148 7789 2150
rect 7813 2148 7869 2150
rect 6826 1128 6882 1184
<< metal3 >>
rect 6637 9890 6703 9893
rect 8226 9890 9026 9920
rect 6637 9888 9026 9890
rect 6637 9832 6642 9888
rect 6698 9832 9026 9888
rect 6637 9830 9026 9832
rect 6637 9827 6703 9830
rect 8226 9800 9026 9830
rect 8017 8802 8083 8805
rect 8226 8802 9026 8832
rect 8017 8800 9026 8802
rect 8017 8744 8022 8800
rect 8078 8744 9026 8800
rect 8017 8742 9026 8744
rect 8017 8739 8083 8742
rect 2457 8736 2773 8737
rect 2457 8672 2463 8736
rect 2527 8672 2543 8736
rect 2607 8672 2623 8736
rect 2687 8672 2703 8736
rect 2767 8672 2773 8736
rect 2457 8671 2773 8672
rect 4159 8736 4475 8737
rect 4159 8672 4165 8736
rect 4229 8672 4245 8736
rect 4309 8672 4325 8736
rect 4389 8672 4405 8736
rect 4469 8672 4475 8736
rect 4159 8671 4475 8672
rect 5861 8736 6177 8737
rect 5861 8672 5867 8736
rect 5931 8672 5947 8736
rect 6011 8672 6027 8736
rect 6091 8672 6107 8736
rect 6171 8672 6177 8736
rect 5861 8671 6177 8672
rect 7563 8736 7879 8737
rect 7563 8672 7569 8736
rect 7633 8672 7649 8736
rect 7713 8672 7729 8736
rect 7793 8672 7809 8736
rect 7873 8672 7879 8736
rect 8226 8712 9026 8742
rect 7563 8671 7879 8672
rect 1797 8192 2113 8193
rect 1797 8128 1803 8192
rect 1867 8128 1883 8192
rect 1947 8128 1963 8192
rect 2027 8128 2043 8192
rect 2107 8128 2113 8192
rect 1797 8127 2113 8128
rect 3499 8192 3815 8193
rect 3499 8128 3505 8192
rect 3569 8128 3585 8192
rect 3649 8128 3665 8192
rect 3729 8128 3745 8192
rect 3809 8128 3815 8192
rect 3499 8127 3815 8128
rect 5201 8192 5517 8193
rect 5201 8128 5207 8192
rect 5271 8128 5287 8192
rect 5351 8128 5367 8192
rect 5431 8128 5447 8192
rect 5511 8128 5517 8192
rect 5201 8127 5517 8128
rect 6903 8192 7219 8193
rect 6903 8128 6909 8192
rect 6973 8128 6989 8192
rect 7053 8128 7069 8192
rect 7133 8128 7149 8192
rect 7213 8128 7219 8192
rect 6903 8127 7219 8128
rect 8017 7714 8083 7717
rect 8226 7714 9026 7744
rect 8017 7712 9026 7714
rect 8017 7656 8022 7712
rect 8078 7656 9026 7712
rect 8017 7654 9026 7656
rect 8017 7651 8083 7654
rect 2457 7648 2773 7649
rect 2457 7584 2463 7648
rect 2527 7584 2543 7648
rect 2607 7584 2623 7648
rect 2687 7584 2703 7648
rect 2767 7584 2773 7648
rect 2457 7583 2773 7584
rect 4159 7648 4475 7649
rect 4159 7584 4165 7648
rect 4229 7584 4245 7648
rect 4309 7584 4325 7648
rect 4389 7584 4405 7648
rect 4469 7584 4475 7648
rect 4159 7583 4475 7584
rect 5861 7648 6177 7649
rect 5861 7584 5867 7648
rect 5931 7584 5947 7648
rect 6011 7584 6027 7648
rect 6091 7584 6107 7648
rect 6171 7584 6177 7648
rect 5861 7583 6177 7584
rect 7563 7648 7879 7649
rect 7563 7584 7569 7648
rect 7633 7584 7649 7648
rect 7713 7584 7729 7648
rect 7793 7584 7809 7648
rect 7873 7584 7879 7648
rect 8226 7624 9026 7654
rect 7563 7583 7879 7584
rect 4429 7442 4495 7445
rect 5257 7442 5323 7445
rect 4429 7440 5323 7442
rect 4429 7384 4434 7440
rect 4490 7384 5262 7440
rect 5318 7384 5323 7440
rect 4429 7382 5323 7384
rect 4429 7379 4495 7382
rect 5257 7379 5323 7382
rect 1797 7104 2113 7105
rect 1797 7040 1803 7104
rect 1867 7040 1883 7104
rect 1947 7040 1963 7104
rect 2027 7040 2043 7104
rect 2107 7040 2113 7104
rect 1797 7039 2113 7040
rect 3499 7104 3815 7105
rect 3499 7040 3505 7104
rect 3569 7040 3585 7104
rect 3649 7040 3665 7104
rect 3729 7040 3745 7104
rect 3809 7040 3815 7104
rect 3499 7039 3815 7040
rect 5201 7104 5517 7105
rect 5201 7040 5207 7104
rect 5271 7040 5287 7104
rect 5351 7040 5367 7104
rect 5431 7040 5447 7104
rect 5511 7040 5517 7104
rect 5201 7039 5517 7040
rect 6903 7104 7219 7105
rect 6903 7040 6909 7104
rect 6973 7040 6989 7104
rect 7053 7040 7069 7104
rect 7133 7040 7149 7104
rect 7213 7040 7219 7104
rect 6903 7039 7219 7040
rect 8017 6626 8083 6629
rect 8226 6626 9026 6656
rect 8017 6624 9026 6626
rect 8017 6568 8022 6624
rect 8078 6568 9026 6624
rect 8017 6566 9026 6568
rect 8017 6563 8083 6566
rect 2457 6560 2773 6561
rect 2457 6496 2463 6560
rect 2527 6496 2543 6560
rect 2607 6496 2623 6560
rect 2687 6496 2703 6560
rect 2767 6496 2773 6560
rect 2457 6495 2773 6496
rect 4159 6560 4475 6561
rect 4159 6496 4165 6560
rect 4229 6496 4245 6560
rect 4309 6496 4325 6560
rect 4389 6496 4405 6560
rect 4469 6496 4475 6560
rect 4159 6495 4475 6496
rect 5861 6560 6177 6561
rect 5861 6496 5867 6560
rect 5931 6496 5947 6560
rect 6011 6496 6027 6560
rect 6091 6496 6107 6560
rect 6171 6496 6177 6560
rect 5861 6495 6177 6496
rect 7563 6560 7879 6561
rect 7563 6496 7569 6560
rect 7633 6496 7649 6560
rect 7713 6496 7729 6560
rect 7793 6496 7809 6560
rect 7873 6496 7879 6560
rect 8226 6536 9026 6566
rect 7563 6495 7879 6496
rect 1797 6016 2113 6017
rect 1797 5952 1803 6016
rect 1867 5952 1883 6016
rect 1947 5952 1963 6016
rect 2027 5952 2043 6016
rect 2107 5952 2113 6016
rect 1797 5951 2113 5952
rect 3499 6016 3815 6017
rect 3499 5952 3505 6016
rect 3569 5952 3585 6016
rect 3649 5952 3665 6016
rect 3729 5952 3745 6016
rect 3809 5952 3815 6016
rect 3499 5951 3815 5952
rect 5201 6016 5517 6017
rect 5201 5952 5207 6016
rect 5271 5952 5287 6016
rect 5351 5952 5367 6016
rect 5431 5952 5447 6016
rect 5511 5952 5517 6016
rect 5201 5951 5517 5952
rect 6903 6016 7219 6017
rect 6903 5952 6909 6016
rect 6973 5952 6989 6016
rect 7053 5952 7069 6016
rect 7133 5952 7149 6016
rect 7213 5952 7219 6016
rect 6903 5951 7219 5952
rect 8017 5538 8083 5541
rect 8226 5538 9026 5568
rect 8017 5536 9026 5538
rect 8017 5480 8022 5536
rect 8078 5480 9026 5536
rect 8017 5478 9026 5480
rect 8017 5475 8083 5478
rect 2457 5472 2773 5473
rect 2457 5408 2463 5472
rect 2527 5408 2543 5472
rect 2607 5408 2623 5472
rect 2687 5408 2703 5472
rect 2767 5408 2773 5472
rect 2457 5407 2773 5408
rect 4159 5472 4475 5473
rect 4159 5408 4165 5472
rect 4229 5408 4245 5472
rect 4309 5408 4325 5472
rect 4389 5408 4405 5472
rect 4469 5408 4475 5472
rect 4159 5407 4475 5408
rect 5861 5472 6177 5473
rect 5861 5408 5867 5472
rect 5931 5408 5947 5472
rect 6011 5408 6027 5472
rect 6091 5408 6107 5472
rect 6171 5408 6177 5472
rect 5861 5407 6177 5408
rect 7563 5472 7879 5473
rect 7563 5408 7569 5472
rect 7633 5408 7649 5472
rect 7713 5408 7729 5472
rect 7793 5408 7809 5472
rect 7873 5408 7879 5472
rect 8226 5448 9026 5478
rect 7563 5407 7879 5408
rect 1797 4928 2113 4929
rect 1797 4864 1803 4928
rect 1867 4864 1883 4928
rect 1947 4864 1963 4928
rect 2027 4864 2043 4928
rect 2107 4864 2113 4928
rect 1797 4863 2113 4864
rect 3499 4928 3815 4929
rect 3499 4864 3505 4928
rect 3569 4864 3585 4928
rect 3649 4864 3665 4928
rect 3729 4864 3745 4928
rect 3809 4864 3815 4928
rect 3499 4863 3815 4864
rect 5201 4928 5517 4929
rect 5201 4864 5207 4928
rect 5271 4864 5287 4928
rect 5351 4864 5367 4928
rect 5431 4864 5447 4928
rect 5511 4864 5517 4928
rect 5201 4863 5517 4864
rect 6903 4928 7219 4929
rect 6903 4864 6909 4928
rect 6973 4864 6989 4928
rect 7053 4864 7069 4928
rect 7133 4864 7149 4928
rect 7213 4864 7219 4928
rect 6903 4863 7219 4864
rect 8017 4450 8083 4453
rect 8226 4450 9026 4480
rect 8017 4448 9026 4450
rect 8017 4392 8022 4448
rect 8078 4392 9026 4448
rect 8017 4390 9026 4392
rect 8017 4387 8083 4390
rect 2457 4384 2773 4385
rect 2457 4320 2463 4384
rect 2527 4320 2543 4384
rect 2607 4320 2623 4384
rect 2687 4320 2703 4384
rect 2767 4320 2773 4384
rect 2457 4319 2773 4320
rect 4159 4384 4475 4385
rect 4159 4320 4165 4384
rect 4229 4320 4245 4384
rect 4309 4320 4325 4384
rect 4389 4320 4405 4384
rect 4469 4320 4475 4384
rect 4159 4319 4475 4320
rect 5861 4384 6177 4385
rect 5861 4320 5867 4384
rect 5931 4320 5947 4384
rect 6011 4320 6027 4384
rect 6091 4320 6107 4384
rect 6171 4320 6177 4384
rect 5861 4319 6177 4320
rect 7563 4384 7879 4385
rect 7563 4320 7569 4384
rect 7633 4320 7649 4384
rect 7713 4320 7729 4384
rect 7793 4320 7809 4384
rect 7873 4320 7879 4384
rect 8226 4360 9026 4390
rect 7563 4319 7879 4320
rect 4429 4178 4495 4181
rect 5625 4178 5691 4181
rect 4429 4176 5691 4178
rect 4429 4120 4434 4176
rect 4490 4120 5630 4176
rect 5686 4120 5691 4176
rect 4429 4118 5691 4120
rect 4429 4115 4495 4118
rect 5625 4115 5691 4118
rect 1797 3840 2113 3841
rect 1797 3776 1803 3840
rect 1867 3776 1883 3840
rect 1947 3776 1963 3840
rect 2027 3776 2043 3840
rect 2107 3776 2113 3840
rect 1797 3775 2113 3776
rect 3499 3840 3815 3841
rect 3499 3776 3505 3840
rect 3569 3776 3585 3840
rect 3649 3776 3665 3840
rect 3729 3776 3745 3840
rect 3809 3776 3815 3840
rect 3499 3775 3815 3776
rect 5201 3840 5517 3841
rect 5201 3776 5207 3840
rect 5271 3776 5287 3840
rect 5351 3776 5367 3840
rect 5431 3776 5447 3840
rect 5511 3776 5517 3840
rect 5201 3775 5517 3776
rect 6903 3840 7219 3841
rect 6903 3776 6909 3840
rect 6973 3776 6989 3840
rect 7053 3776 7069 3840
rect 7133 3776 7149 3840
rect 7213 3776 7219 3840
rect 6903 3775 7219 3776
rect 8017 3362 8083 3365
rect 8226 3362 9026 3392
rect 8017 3360 9026 3362
rect 8017 3304 8022 3360
rect 8078 3304 9026 3360
rect 8017 3302 9026 3304
rect 8017 3299 8083 3302
rect 2457 3296 2773 3297
rect 2457 3232 2463 3296
rect 2527 3232 2543 3296
rect 2607 3232 2623 3296
rect 2687 3232 2703 3296
rect 2767 3232 2773 3296
rect 2457 3231 2773 3232
rect 4159 3296 4475 3297
rect 4159 3232 4165 3296
rect 4229 3232 4245 3296
rect 4309 3232 4325 3296
rect 4389 3232 4405 3296
rect 4469 3232 4475 3296
rect 4159 3231 4475 3232
rect 5861 3296 6177 3297
rect 5861 3232 5867 3296
rect 5931 3232 5947 3296
rect 6011 3232 6027 3296
rect 6091 3232 6107 3296
rect 6171 3232 6177 3296
rect 5861 3231 6177 3232
rect 7563 3296 7879 3297
rect 7563 3232 7569 3296
rect 7633 3232 7649 3296
rect 7713 3232 7729 3296
rect 7793 3232 7809 3296
rect 7873 3232 7879 3296
rect 8226 3272 9026 3302
rect 7563 3231 7879 3232
rect 1797 2752 2113 2753
rect 1797 2688 1803 2752
rect 1867 2688 1883 2752
rect 1947 2688 1963 2752
rect 2027 2688 2043 2752
rect 2107 2688 2113 2752
rect 1797 2687 2113 2688
rect 3499 2752 3815 2753
rect 3499 2688 3505 2752
rect 3569 2688 3585 2752
rect 3649 2688 3665 2752
rect 3729 2688 3745 2752
rect 3809 2688 3815 2752
rect 3499 2687 3815 2688
rect 5201 2752 5517 2753
rect 5201 2688 5207 2752
rect 5271 2688 5287 2752
rect 5351 2688 5367 2752
rect 5431 2688 5447 2752
rect 5511 2688 5517 2752
rect 5201 2687 5517 2688
rect 6903 2752 7219 2753
rect 6903 2688 6909 2752
rect 6973 2688 6989 2752
rect 7053 2688 7069 2752
rect 7133 2688 7149 2752
rect 7213 2688 7219 2752
rect 6903 2687 7219 2688
rect 8017 2274 8083 2277
rect 8226 2274 9026 2304
rect 8017 2272 9026 2274
rect 8017 2216 8022 2272
rect 8078 2216 9026 2272
rect 8017 2214 9026 2216
rect 8017 2211 8083 2214
rect 2457 2208 2773 2209
rect 2457 2144 2463 2208
rect 2527 2144 2543 2208
rect 2607 2144 2623 2208
rect 2687 2144 2703 2208
rect 2767 2144 2773 2208
rect 2457 2143 2773 2144
rect 4159 2208 4475 2209
rect 4159 2144 4165 2208
rect 4229 2144 4245 2208
rect 4309 2144 4325 2208
rect 4389 2144 4405 2208
rect 4469 2144 4475 2208
rect 4159 2143 4475 2144
rect 5861 2208 6177 2209
rect 5861 2144 5867 2208
rect 5931 2144 5947 2208
rect 6011 2144 6027 2208
rect 6091 2144 6107 2208
rect 6171 2144 6177 2208
rect 5861 2143 6177 2144
rect 7563 2208 7879 2209
rect 7563 2144 7569 2208
rect 7633 2144 7649 2208
rect 7713 2144 7729 2208
rect 7793 2144 7809 2208
rect 7873 2144 7879 2208
rect 8226 2184 9026 2214
rect 7563 2143 7879 2144
rect 6821 1186 6887 1189
rect 8226 1186 9026 1216
rect 6821 1184 9026 1186
rect 6821 1128 6826 1184
rect 6882 1128 9026 1184
rect 6821 1126 9026 1128
rect 6821 1123 6887 1126
rect 8226 1096 9026 1126
<< via3 >>
rect 2463 8732 2527 8736
rect 2463 8676 2467 8732
rect 2467 8676 2523 8732
rect 2523 8676 2527 8732
rect 2463 8672 2527 8676
rect 2543 8732 2607 8736
rect 2543 8676 2547 8732
rect 2547 8676 2603 8732
rect 2603 8676 2607 8732
rect 2543 8672 2607 8676
rect 2623 8732 2687 8736
rect 2623 8676 2627 8732
rect 2627 8676 2683 8732
rect 2683 8676 2687 8732
rect 2623 8672 2687 8676
rect 2703 8732 2767 8736
rect 2703 8676 2707 8732
rect 2707 8676 2763 8732
rect 2763 8676 2767 8732
rect 2703 8672 2767 8676
rect 4165 8732 4229 8736
rect 4165 8676 4169 8732
rect 4169 8676 4225 8732
rect 4225 8676 4229 8732
rect 4165 8672 4229 8676
rect 4245 8732 4309 8736
rect 4245 8676 4249 8732
rect 4249 8676 4305 8732
rect 4305 8676 4309 8732
rect 4245 8672 4309 8676
rect 4325 8732 4389 8736
rect 4325 8676 4329 8732
rect 4329 8676 4385 8732
rect 4385 8676 4389 8732
rect 4325 8672 4389 8676
rect 4405 8732 4469 8736
rect 4405 8676 4409 8732
rect 4409 8676 4465 8732
rect 4465 8676 4469 8732
rect 4405 8672 4469 8676
rect 5867 8732 5931 8736
rect 5867 8676 5871 8732
rect 5871 8676 5927 8732
rect 5927 8676 5931 8732
rect 5867 8672 5931 8676
rect 5947 8732 6011 8736
rect 5947 8676 5951 8732
rect 5951 8676 6007 8732
rect 6007 8676 6011 8732
rect 5947 8672 6011 8676
rect 6027 8732 6091 8736
rect 6027 8676 6031 8732
rect 6031 8676 6087 8732
rect 6087 8676 6091 8732
rect 6027 8672 6091 8676
rect 6107 8732 6171 8736
rect 6107 8676 6111 8732
rect 6111 8676 6167 8732
rect 6167 8676 6171 8732
rect 6107 8672 6171 8676
rect 7569 8732 7633 8736
rect 7569 8676 7573 8732
rect 7573 8676 7629 8732
rect 7629 8676 7633 8732
rect 7569 8672 7633 8676
rect 7649 8732 7713 8736
rect 7649 8676 7653 8732
rect 7653 8676 7709 8732
rect 7709 8676 7713 8732
rect 7649 8672 7713 8676
rect 7729 8732 7793 8736
rect 7729 8676 7733 8732
rect 7733 8676 7789 8732
rect 7789 8676 7793 8732
rect 7729 8672 7793 8676
rect 7809 8732 7873 8736
rect 7809 8676 7813 8732
rect 7813 8676 7869 8732
rect 7869 8676 7873 8732
rect 7809 8672 7873 8676
rect 1803 8188 1867 8192
rect 1803 8132 1807 8188
rect 1807 8132 1863 8188
rect 1863 8132 1867 8188
rect 1803 8128 1867 8132
rect 1883 8188 1947 8192
rect 1883 8132 1887 8188
rect 1887 8132 1943 8188
rect 1943 8132 1947 8188
rect 1883 8128 1947 8132
rect 1963 8188 2027 8192
rect 1963 8132 1967 8188
rect 1967 8132 2023 8188
rect 2023 8132 2027 8188
rect 1963 8128 2027 8132
rect 2043 8188 2107 8192
rect 2043 8132 2047 8188
rect 2047 8132 2103 8188
rect 2103 8132 2107 8188
rect 2043 8128 2107 8132
rect 3505 8188 3569 8192
rect 3505 8132 3509 8188
rect 3509 8132 3565 8188
rect 3565 8132 3569 8188
rect 3505 8128 3569 8132
rect 3585 8188 3649 8192
rect 3585 8132 3589 8188
rect 3589 8132 3645 8188
rect 3645 8132 3649 8188
rect 3585 8128 3649 8132
rect 3665 8188 3729 8192
rect 3665 8132 3669 8188
rect 3669 8132 3725 8188
rect 3725 8132 3729 8188
rect 3665 8128 3729 8132
rect 3745 8188 3809 8192
rect 3745 8132 3749 8188
rect 3749 8132 3805 8188
rect 3805 8132 3809 8188
rect 3745 8128 3809 8132
rect 5207 8188 5271 8192
rect 5207 8132 5211 8188
rect 5211 8132 5267 8188
rect 5267 8132 5271 8188
rect 5207 8128 5271 8132
rect 5287 8188 5351 8192
rect 5287 8132 5291 8188
rect 5291 8132 5347 8188
rect 5347 8132 5351 8188
rect 5287 8128 5351 8132
rect 5367 8188 5431 8192
rect 5367 8132 5371 8188
rect 5371 8132 5427 8188
rect 5427 8132 5431 8188
rect 5367 8128 5431 8132
rect 5447 8188 5511 8192
rect 5447 8132 5451 8188
rect 5451 8132 5507 8188
rect 5507 8132 5511 8188
rect 5447 8128 5511 8132
rect 6909 8188 6973 8192
rect 6909 8132 6913 8188
rect 6913 8132 6969 8188
rect 6969 8132 6973 8188
rect 6909 8128 6973 8132
rect 6989 8188 7053 8192
rect 6989 8132 6993 8188
rect 6993 8132 7049 8188
rect 7049 8132 7053 8188
rect 6989 8128 7053 8132
rect 7069 8188 7133 8192
rect 7069 8132 7073 8188
rect 7073 8132 7129 8188
rect 7129 8132 7133 8188
rect 7069 8128 7133 8132
rect 7149 8188 7213 8192
rect 7149 8132 7153 8188
rect 7153 8132 7209 8188
rect 7209 8132 7213 8188
rect 7149 8128 7213 8132
rect 2463 7644 2527 7648
rect 2463 7588 2467 7644
rect 2467 7588 2523 7644
rect 2523 7588 2527 7644
rect 2463 7584 2527 7588
rect 2543 7644 2607 7648
rect 2543 7588 2547 7644
rect 2547 7588 2603 7644
rect 2603 7588 2607 7644
rect 2543 7584 2607 7588
rect 2623 7644 2687 7648
rect 2623 7588 2627 7644
rect 2627 7588 2683 7644
rect 2683 7588 2687 7644
rect 2623 7584 2687 7588
rect 2703 7644 2767 7648
rect 2703 7588 2707 7644
rect 2707 7588 2763 7644
rect 2763 7588 2767 7644
rect 2703 7584 2767 7588
rect 4165 7644 4229 7648
rect 4165 7588 4169 7644
rect 4169 7588 4225 7644
rect 4225 7588 4229 7644
rect 4165 7584 4229 7588
rect 4245 7644 4309 7648
rect 4245 7588 4249 7644
rect 4249 7588 4305 7644
rect 4305 7588 4309 7644
rect 4245 7584 4309 7588
rect 4325 7644 4389 7648
rect 4325 7588 4329 7644
rect 4329 7588 4385 7644
rect 4385 7588 4389 7644
rect 4325 7584 4389 7588
rect 4405 7644 4469 7648
rect 4405 7588 4409 7644
rect 4409 7588 4465 7644
rect 4465 7588 4469 7644
rect 4405 7584 4469 7588
rect 5867 7644 5931 7648
rect 5867 7588 5871 7644
rect 5871 7588 5927 7644
rect 5927 7588 5931 7644
rect 5867 7584 5931 7588
rect 5947 7644 6011 7648
rect 5947 7588 5951 7644
rect 5951 7588 6007 7644
rect 6007 7588 6011 7644
rect 5947 7584 6011 7588
rect 6027 7644 6091 7648
rect 6027 7588 6031 7644
rect 6031 7588 6087 7644
rect 6087 7588 6091 7644
rect 6027 7584 6091 7588
rect 6107 7644 6171 7648
rect 6107 7588 6111 7644
rect 6111 7588 6167 7644
rect 6167 7588 6171 7644
rect 6107 7584 6171 7588
rect 7569 7644 7633 7648
rect 7569 7588 7573 7644
rect 7573 7588 7629 7644
rect 7629 7588 7633 7644
rect 7569 7584 7633 7588
rect 7649 7644 7713 7648
rect 7649 7588 7653 7644
rect 7653 7588 7709 7644
rect 7709 7588 7713 7644
rect 7649 7584 7713 7588
rect 7729 7644 7793 7648
rect 7729 7588 7733 7644
rect 7733 7588 7789 7644
rect 7789 7588 7793 7644
rect 7729 7584 7793 7588
rect 7809 7644 7873 7648
rect 7809 7588 7813 7644
rect 7813 7588 7869 7644
rect 7869 7588 7873 7644
rect 7809 7584 7873 7588
rect 1803 7100 1867 7104
rect 1803 7044 1807 7100
rect 1807 7044 1863 7100
rect 1863 7044 1867 7100
rect 1803 7040 1867 7044
rect 1883 7100 1947 7104
rect 1883 7044 1887 7100
rect 1887 7044 1943 7100
rect 1943 7044 1947 7100
rect 1883 7040 1947 7044
rect 1963 7100 2027 7104
rect 1963 7044 1967 7100
rect 1967 7044 2023 7100
rect 2023 7044 2027 7100
rect 1963 7040 2027 7044
rect 2043 7100 2107 7104
rect 2043 7044 2047 7100
rect 2047 7044 2103 7100
rect 2103 7044 2107 7100
rect 2043 7040 2107 7044
rect 3505 7100 3569 7104
rect 3505 7044 3509 7100
rect 3509 7044 3565 7100
rect 3565 7044 3569 7100
rect 3505 7040 3569 7044
rect 3585 7100 3649 7104
rect 3585 7044 3589 7100
rect 3589 7044 3645 7100
rect 3645 7044 3649 7100
rect 3585 7040 3649 7044
rect 3665 7100 3729 7104
rect 3665 7044 3669 7100
rect 3669 7044 3725 7100
rect 3725 7044 3729 7100
rect 3665 7040 3729 7044
rect 3745 7100 3809 7104
rect 3745 7044 3749 7100
rect 3749 7044 3805 7100
rect 3805 7044 3809 7100
rect 3745 7040 3809 7044
rect 5207 7100 5271 7104
rect 5207 7044 5211 7100
rect 5211 7044 5267 7100
rect 5267 7044 5271 7100
rect 5207 7040 5271 7044
rect 5287 7100 5351 7104
rect 5287 7044 5291 7100
rect 5291 7044 5347 7100
rect 5347 7044 5351 7100
rect 5287 7040 5351 7044
rect 5367 7100 5431 7104
rect 5367 7044 5371 7100
rect 5371 7044 5427 7100
rect 5427 7044 5431 7100
rect 5367 7040 5431 7044
rect 5447 7100 5511 7104
rect 5447 7044 5451 7100
rect 5451 7044 5507 7100
rect 5507 7044 5511 7100
rect 5447 7040 5511 7044
rect 6909 7100 6973 7104
rect 6909 7044 6913 7100
rect 6913 7044 6969 7100
rect 6969 7044 6973 7100
rect 6909 7040 6973 7044
rect 6989 7100 7053 7104
rect 6989 7044 6993 7100
rect 6993 7044 7049 7100
rect 7049 7044 7053 7100
rect 6989 7040 7053 7044
rect 7069 7100 7133 7104
rect 7069 7044 7073 7100
rect 7073 7044 7129 7100
rect 7129 7044 7133 7100
rect 7069 7040 7133 7044
rect 7149 7100 7213 7104
rect 7149 7044 7153 7100
rect 7153 7044 7209 7100
rect 7209 7044 7213 7100
rect 7149 7040 7213 7044
rect 2463 6556 2527 6560
rect 2463 6500 2467 6556
rect 2467 6500 2523 6556
rect 2523 6500 2527 6556
rect 2463 6496 2527 6500
rect 2543 6556 2607 6560
rect 2543 6500 2547 6556
rect 2547 6500 2603 6556
rect 2603 6500 2607 6556
rect 2543 6496 2607 6500
rect 2623 6556 2687 6560
rect 2623 6500 2627 6556
rect 2627 6500 2683 6556
rect 2683 6500 2687 6556
rect 2623 6496 2687 6500
rect 2703 6556 2767 6560
rect 2703 6500 2707 6556
rect 2707 6500 2763 6556
rect 2763 6500 2767 6556
rect 2703 6496 2767 6500
rect 4165 6556 4229 6560
rect 4165 6500 4169 6556
rect 4169 6500 4225 6556
rect 4225 6500 4229 6556
rect 4165 6496 4229 6500
rect 4245 6556 4309 6560
rect 4245 6500 4249 6556
rect 4249 6500 4305 6556
rect 4305 6500 4309 6556
rect 4245 6496 4309 6500
rect 4325 6556 4389 6560
rect 4325 6500 4329 6556
rect 4329 6500 4385 6556
rect 4385 6500 4389 6556
rect 4325 6496 4389 6500
rect 4405 6556 4469 6560
rect 4405 6500 4409 6556
rect 4409 6500 4465 6556
rect 4465 6500 4469 6556
rect 4405 6496 4469 6500
rect 5867 6556 5931 6560
rect 5867 6500 5871 6556
rect 5871 6500 5927 6556
rect 5927 6500 5931 6556
rect 5867 6496 5931 6500
rect 5947 6556 6011 6560
rect 5947 6500 5951 6556
rect 5951 6500 6007 6556
rect 6007 6500 6011 6556
rect 5947 6496 6011 6500
rect 6027 6556 6091 6560
rect 6027 6500 6031 6556
rect 6031 6500 6087 6556
rect 6087 6500 6091 6556
rect 6027 6496 6091 6500
rect 6107 6556 6171 6560
rect 6107 6500 6111 6556
rect 6111 6500 6167 6556
rect 6167 6500 6171 6556
rect 6107 6496 6171 6500
rect 7569 6556 7633 6560
rect 7569 6500 7573 6556
rect 7573 6500 7629 6556
rect 7629 6500 7633 6556
rect 7569 6496 7633 6500
rect 7649 6556 7713 6560
rect 7649 6500 7653 6556
rect 7653 6500 7709 6556
rect 7709 6500 7713 6556
rect 7649 6496 7713 6500
rect 7729 6556 7793 6560
rect 7729 6500 7733 6556
rect 7733 6500 7789 6556
rect 7789 6500 7793 6556
rect 7729 6496 7793 6500
rect 7809 6556 7873 6560
rect 7809 6500 7813 6556
rect 7813 6500 7869 6556
rect 7869 6500 7873 6556
rect 7809 6496 7873 6500
rect 1803 6012 1867 6016
rect 1803 5956 1807 6012
rect 1807 5956 1863 6012
rect 1863 5956 1867 6012
rect 1803 5952 1867 5956
rect 1883 6012 1947 6016
rect 1883 5956 1887 6012
rect 1887 5956 1943 6012
rect 1943 5956 1947 6012
rect 1883 5952 1947 5956
rect 1963 6012 2027 6016
rect 1963 5956 1967 6012
rect 1967 5956 2023 6012
rect 2023 5956 2027 6012
rect 1963 5952 2027 5956
rect 2043 6012 2107 6016
rect 2043 5956 2047 6012
rect 2047 5956 2103 6012
rect 2103 5956 2107 6012
rect 2043 5952 2107 5956
rect 3505 6012 3569 6016
rect 3505 5956 3509 6012
rect 3509 5956 3565 6012
rect 3565 5956 3569 6012
rect 3505 5952 3569 5956
rect 3585 6012 3649 6016
rect 3585 5956 3589 6012
rect 3589 5956 3645 6012
rect 3645 5956 3649 6012
rect 3585 5952 3649 5956
rect 3665 6012 3729 6016
rect 3665 5956 3669 6012
rect 3669 5956 3725 6012
rect 3725 5956 3729 6012
rect 3665 5952 3729 5956
rect 3745 6012 3809 6016
rect 3745 5956 3749 6012
rect 3749 5956 3805 6012
rect 3805 5956 3809 6012
rect 3745 5952 3809 5956
rect 5207 6012 5271 6016
rect 5207 5956 5211 6012
rect 5211 5956 5267 6012
rect 5267 5956 5271 6012
rect 5207 5952 5271 5956
rect 5287 6012 5351 6016
rect 5287 5956 5291 6012
rect 5291 5956 5347 6012
rect 5347 5956 5351 6012
rect 5287 5952 5351 5956
rect 5367 6012 5431 6016
rect 5367 5956 5371 6012
rect 5371 5956 5427 6012
rect 5427 5956 5431 6012
rect 5367 5952 5431 5956
rect 5447 6012 5511 6016
rect 5447 5956 5451 6012
rect 5451 5956 5507 6012
rect 5507 5956 5511 6012
rect 5447 5952 5511 5956
rect 6909 6012 6973 6016
rect 6909 5956 6913 6012
rect 6913 5956 6969 6012
rect 6969 5956 6973 6012
rect 6909 5952 6973 5956
rect 6989 6012 7053 6016
rect 6989 5956 6993 6012
rect 6993 5956 7049 6012
rect 7049 5956 7053 6012
rect 6989 5952 7053 5956
rect 7069 6012 7133 6016
rect 7069 5956 7073 6012
rect 7073 5956 7129 6012
rect 7129 5956 7133 6012
rect 7069 5952 7133 5956
rect 7149 6012 7213 6016
rect 7149 5956 7153 6012
rect 7153 5956 7209 6012
rect 7209 5956 7213 6012
rect 7149 5952 7213 5956
rect 2463 5468 2527 5472
rect 2463 5412 2467 5468
rect 2467 5412 2523 5468
rect 2523 5412 2527 5468
rect 2463 5408 2527 5412
rect 2543 5468 2607 5472
rect 2543 5412 2547 5468
rect 2547 5412 2603 5468
rect 2603 5412 2607 5468
rect 2543 5408 2607 5412
rect 2623 5468 2687 5472
rect 2623 5412 2627 5468
rect 2627 5412 2683 5468
rect 2683 5412 2687 5468
rect 2623 5408 2687 5412
rect 2703 5468 2767 5472
rect 2703 5412 2707 5468
rect 2707 5412 2763 5468
rect 2763 5412 2767 5468
rect 2703 5408 2767 5412
rect 4165 5468 4229 5472
rect 4165 5412 4169 5468
rect 4169 5412 4225 5468
rect 4225 5412 4229 5468
rect 4165 5408 4229 5412
rect 4245 5468 4309 5472
rect 4245 5412 4249 5468
rect 4249 5412 4305 5468
rect 4305 5412 4309 5468
rect 4245 5408 4309 5412
rect 4325 5468 4389 5472
rect 4325 5412 4329 5468
rect 4329 5412 4385 5468
rect 4385 5412 4389 5468
rect 4325 5408 4389 5412
rect 4405 5468 4469 5472
rect 4405 5412 4409 5468
rect 4409 5412 4465 5468
rect 4465 5412 4469 5468
rect 4405 5408 4469 5412
rect 5867 5468 5931 5472
rect 5867 5412 5871 5468
rect 5871 5412 5927 5468
rect 5927 5412 5931 5468
rect 5867 5408 5931 5412
rect 5947 5468 6011 5472
rect 5947 5412 5951 5468
rect 5951 5412 6007 5468
rect 6007 5412 6011 5468
rect 5947 5408 6011 5412
rect 6027 5468 6091 5472
rect 6027 5412 6031 5468
rect 6031 5412 6087 5468
rect 6087 5412 6091 5468
rect 6027 5408 6091 5412
rect 6107 5468 6171 5472
rect 6107 5412 6111 5468
rect 6111 5412 6167 5468
rect 6167 5412 6171 5468
rect 6107 5408 6171 5412
rect 7569 5468 7633 5472
rect 7569 5412 7573 5468
rect 7573 5412 7629 5468
rect 7629 5412 7633 5468
rect 7569 5408 7633 5412
rect 7649 5468 7713 5472
rect 7649 5412 7653 5468
rect 7653 5412 7709 5468
rect 7709 5412 7713 5468
rect 7649 5408 7713 5412
rect 7729 5468 7793 5472
rect 7729 5412 7733 5468
rect 7733 5412 7789 5468
rect 7789 5412 7793 5468
rect 7729 5408 7793 5412
rect 7809 5468 7873 5472
rect 7809 5412 7813 5468
rect 7813 5412 7869 5468
rect 7869 5412 7873 5468
rect 7809 5408 7873 5412
rect 1803 4924 1867 4928
rect 1803 4868 1807 4924
rect 1807 4868 1863 4924
rect 1863 4868 1867 4924
rect 1803 4864 1867 4868
rect 1883 4924 1947 4928
rect 1883 4868 1887 4924
rect 1887 4868 1943 4924
rect 1943 4868 1947 4924
rect 1883 4864 1947 4868
rect 1963 4924 2027 4928
rect 1963 4868 1967 4924
rect 1967 4868 2023 4924
rect 2023 4868 2027 4924
rect 1963 4864 2027 4868
rect 2043 4924 2107 4928
rect 2043 4868 2047 4924
rect 2047 4868 2103 4924
rect 2103 4868 2107 4924
rect 2043 4864 2107 4868
rect 3505 4924 3569 4928
rect 3505 4868 3509 4924
rect 3509 4868 3565 4924
rect 3565 4868 3569 4924
rect 3505 4864 3569 4868
rect 3585 4924 3649 4928
rect 3585 4868 3589 4924
rect 3589 4868 3645 4924
rect 3645 4868 3649 4924
rect 3585 4864 3649 4868
rect 3665 4924 3729 4928
rect 3665 4868 3669 4924
rect 3669 4868 3725 4924
rect 3725 4868 3729 4924
rect 3665 4864 3729 4868
rect 3745 4924 3809 4928
rect 3745 4868 3749 4924
rect 3749 4868 3805 4924
rect 3805 4868 3809 4924
rect 3745 4864 3809 4868
rect 5207 4924 5271 4928
rect 5207 4868 5211 4924
rect 5211 4868 5267 4924
rect 5267 4868 5271 4924
rect 5207 4864 5271 4868
rect 5287 4924 5351 4928
rect 5287 4868 5291 4924
rect 5291 4868 5347 4924
rect 5347 4868 5351 4924
rect 5287 4864 5351 4868
rect 5367 4924 5431 4928
rect 5367 4868 5371 4924
rect 5371 4868 5427 4924
rect 5427 4868 5431 4924
rect 5367 4864 5431 4868
rect 5447 4924 5511 4928
rect 5447 4868 5451 4924
rect 5451 4868 5507 4924
rect 5507 4868 5511 4924
rect 5447 4864 5511 4868
rect 6909 4924 6973 4928
rect 6909 4868 6913 4924
rect 6913 4868 6969 4924
rect 6969 4868 6973 4924
rect 6909 4864 6973 4868
rect 6989 4924 7053 4928
rect 6989 4868 6993 4924
rect 6993 4868 7049 4924
rect 7049 4868 7053 4924
rect 6989 4864 7053 4868
rect 7069 4924 7133 4928
rect 7069 4868 7073 4924
rect 7073 4868 7129 4924
rect 7129 4868 7133 4924
rect 7069 4864 7133 4868
rect 7149 4924 7213 4928
rect 7149 4868 7153 4924
rect 7153 4868 7209 4924
rect 7209 4868 7213 4924
rect 7149 4864 7213 4868
rect 2463 4380 2527 4384
rect 2463 4324 2467 4380
rect 2467 4324 2523 4380
rect 2523 4324 2527 4380
rect 2463 4320 2527 4324
rect 2543 4380 2607 4384
rect 2543 4324 2547 4380
rect 2547 4324 2603 4380
rect 2603 4324 2607 4380
rect 2543 4320 2607 4324
rect 2623 4380 2687 4384
rect 2623 4324 2627 4380
rect 2627 4324 2683 4380
rect 2683 4324 2687 4380
rect 2623 4320 2687 4324
rect 2703 4380 2767 4384
rect 2703 4324 2707 4380
rect 2707 4324 2763 4380
rect 2763 4324 2767 4380
rect 2703 4320 2767 4324
rect 4165 4380 4229 4384
rect 4165 4324 4169 4380
rect 4169 4324 4225 4380
rect 4225 4324 4229 4380
rect 4165 4320 4229 4324
rect 4245 4380 4309 4384
rect 4245 4324 4249 4380
rect 4249 4324 4305 4380
rect 4305 4324 4309 4380
rect 4245 4320 4309 4324
rect 4325 4380 4389 4384
rect 4325 4324 4329 4380
rect 4329 4324 4385 4380
rect 4385 4324 4389 4380
rect 4325 4320 4389 4324
rect 4405 4380 4469 4384
rect 4405 4324 4409 4380
rect 4409 4324 4465 4380
rect 4465 4324 4469 4380
rect 4405 4320 4469 4324
rect 5867 4380 5931 4384
rect 5867 4324 5871 4380
rect 5871 4324 5927 4380
rect 5927 4324 5931 4380
rect 5867 4320 5931 4324
rect 5947 4380 6011 4384
rect 5947 4324 5951 4380
rect 5951 4324 6007 4380
rect 6007 4324 6011 4380
rect 5947 4320 6011 4324
rect 6027 4380 6091 4384
rect 6027 4324 6031 4380
rect 6031 4324 6087 4380
rect 6087 4324 6091 4380
rect 6027 4320 6091 4324
rect 6107 4380 6171 4384
rect 6107 4324 6111 4380
rect 6111 4324 6167 4380
rect 6167 4324 6171 4380
rect 6107 4320 6171 4324
rect 7569 4380 7633 4384
rect 7569 4324 7573 4380
rect 7573 4324 7629 4380
rect 7629 4324 7633 4380
rect 7569 4320 7633 4324
rect 7649 4380 7713 4384
rect 7649 4324 7653 4380
rect 7653 4324 7709 4380
rect 7709 4324 7713 4380
rect 7649 4320 7713 4324
rect 7729 4380 7793 4384
rect 7729 4324 7733 4380
rect 7733 4324 7789 4380
rect 7789 4324 7793 4380
rect 7729 4320 7793 4324
rect 7809 4380 7873 4384
rect 7809 4324 7813 4380
rect 7813 4324 7869 4380
rect 7869 4324 7873 4380
rect 7809 4320 7873 4324
rect 1803 3836 1867 3840
rect 1803 3780 1807 3836
rect 1807 3780 1863 3836
rect 1863 3780 1867 3836
rect 1803 3776 1867 3780
rect 1883 3836 1947 3840
rect 1883 3780 1887 3836
rect 1887 3780 1943 3836
rect 1943 3780 1947 3836
rect 1883 3776 1947 3780
rect 1963 3836 2027 3840
rect 1963 3780 1967 3836
rect 1967 3780 2023 3836
rect 2023 3780 2027 3836
rect 1963 3776 2027 3780
rect 2043 3836 2107 3840
rect 2043 3780 2047 3836
rect 2047 3780 2103 3836
rect 2103 3780 2107 3836
rect 2043 3776 2107 3780
rect 3505 3836 3569 3840
rect 3505 3780 3509 3836
rect 3509 3780 3565 3836
rect 3565 3780 3569 3836
rect 3505 3776 3569 3780
rect 3585 3836 3649 3840
rect 3585 3780 3589 3836
rect 3589 3780 3645 3836
rect 3645 3780 3649 3836
rect 3585 3776 3649 3780
rect 3665 3836 3729 3840
rect 3665 3780 3669 3836
rect 3669 3780 3725 3836
rect 3725 3780 3729 3836
rect 3665 3776 3729 3780
rect 3745 3836 3809 3840
rect 3745 3780 3749 3836
rect 3749 3780 3805 3836
rect 3805 3780 3809 3836
rect 3745 3776 3809 3780
rect 5207 3836 5271 3840
rect 5207 3780 5211 3836
rect 5211 3780 5267 3836
rect 5267 3780 5271 3836
rect 5207 3776 5271 3780
rect 5287 3836 5351 3840
rect 5287 3780 5291 3836
rect 5291 3780 5347 3836
rect 5347 3780 5351 3836
rect 5287 3776 5351 3780
rect 5367 3836 5431 3840
rect 5367 3780 5371 3836
rect 5371 3780 5427 3836
rect 5427 3780 5431 3836
rect 5367 3776 5431 3780
rect 5447 3836 5511 3840
rect 5447 3780 5451 3836
rect 5451 3780 5507 3836
rect 5507 3780 5511 3836
rect 5447 3776 5511 3780
rect 6909 3836 6973 3840
rect 6909 3780 6913 3836
rect 6913 3780 6969 3836
rect 6969 3780 6973 3836
rect 6909 3776 6973 3780
rect 6989 3836 7053 3840
rect 6989 3780 6993 3836
rect 6993 3780 7049 3836
rect 7049 3780 7053 3836
rect 6989 3776 7053 3780
rect 7069 3836 7133 3840
rect 7069 3780 7073 3836
rect 7073 3780 7129 3836
rect 7129 3780 7133 3836
rect 7069 3776 7133 3780
rect 7149 3836 7213 3840
rect 7149 3780 7153 3836
rect 7153 3780 7209 3836
rect 7209 3780 7213 3836
rect 7149 3776 7213 3780
rect 2463 3292 2527 3296
rect 2463 3236 2467 3292
rect 2467 3236 2523 3292
rect 2523 3236 2527 3292
rect 2463 3232 2527 3236
rect 2543 3292 2607 3296
rect 2543 3236 2547 3292
rect 2547 3236 2603 3292
rect 2603 3236 2607 3292
rect 2543 3232 2607 3236
rect 2623 3292 2687 3296
rect 2623 3236 2627 3292
rect 2627 3236 2683 3292
rect 2683 3236 2687 3292
rect 2623 3232 2687 3236
rect 2703 3292 2767 3296
rect 2703 3236 2707 3292
rect 2707 3236 2763 3292
rect 2763 3236 2767 3292
rect 2703 3232 2767 3236
rect 4165 3292 4229 3296
rect 4165 3236 4169 3292
rect 4169 3236 4225 3292
rect 4225 3236 4229 3292
rect 4165 3232 4229 3236
rect 4245 3292 4309 3296
rect 4245 3236 4249 3292
rect 4249 3236 4305 3292
rect 4305 3236 4309 3292
rect 4245 3232 4309 3236
rect 4325 3292 4389 3296
rect 4325 3236 4329 3292
rect 4329 3236 4385 3292
rect 4385 3236 4389 3292
rect 4325 3232 4389 3236
rect 4405 3292 4469 3296
rect 4405 3236 4409 3292
rect 4409 3236 4465 3292
rect 4465 3236 4469 3292
rect 4405 3232 4469 3236
rect 5867 3292 5931 3296
rect 5867 3236 5871 3292
rect 5871 3236 5927 3292
rect 5927 3236 5931 3292
rect 5867 3232 5931 3236
rect 5947 3292 6011 3296
rect 5947 3236 5951 3292
rect 5951 3236 6007 3292
rect 6007 3236 6011 3292
rect 5947 3232 6011 3236
rect 6027 3292 6091 3296
rect 6027 3236 6031 3292
rect 6031 3236 6087 3292
rect 6087 3236 6091 3292
rect 6027 3232 6091 3236
rect 6107 3292 6171 3296
rect 6107 3236 6111 3292
rect 6111 3236 6167 3292
rect 6167 3236 6171 3292
rect 6107 3232 6171 3236
rect 7569 3292 7633 3296
rect 7569 3236 7573 3292
rect 7573 3236 7629 3292
rect 7629 3236 7633 3292
rect 7569 3232 7633 3236
rect 7649 3292 7713 3296
rect 7649 3236 7653 3292
rect 7653 3236 7709 3292
rect 7709 3236 7713 3292
rect 7649 3232 7713 3236
rect 7729 3292 7793 3296
rect 7729 3236 7733 3292
rect 7733 3236 7789 3292
rect 7789 3236 7793 3292
rect 7729 3232 7793 3236
rect 7809 3292 7873 3296
rect 7809 3236 7813 3292
rect 7813 3236 7869 3292
rect 7869 3236 7873 3292
rect 7809 3232 7873 3236
rect 1803 2748 1867 2752
rect 1803 2692 1807 2748
rect 1807 2692 1863 2748
rect 1863 2692 1867 2748
rect 1803 2688 1867 2692
rect 1883 2748 1947 2752
rect 1883 2692 1887 2748
rect 1887 2692 1943 2748
rect 1943 2692 1947 2748
rect 1883 2688 1947 2692
rect 1963 2748 2027 2752
rect 1963 2692 1967 2748
rect 1967 2692 2023 2748
rect 2023 2692 2027 2748
rect 1963 2688 2027 2692
rect 2043 2748 2107 2752
rect 2043 2692 2047 2748
rect 2047 2692 2103 2748
rect 2103 2692 2107 2748
rect 2043 2688 2107 2692
rect 3505 2748 3569 2752
rect 3505 2692 3509 2748
rect 3509 2692 3565 2748
rect 3565 2692 3569 2748
rect 3505 2688 3569 2692
rect 3585 2748 3649 2752
rect 3585 2692 3589 2748
rect 3589 2692 3645 2748
rect 3645 2692 3649 2748
rect 3585 2688 3649 2692
rect 3665 2748 3729 2752
rect 3665 2692 3669 2748
rect 3669 2692 3725 2748
rect 3725 2692 3729 2748
rect 3665 2688 3729 2692
rect 3745 2748 3809 2752
rect 3745 2692 3749 2748
rect 3749 2692 3805 2748
rect 3805 2692 3809 2748
rect 3745 2688 3809 2692
rect 5207 2748 5271 2752
rect 5207 2692 5211 2748
rect 5211 2692 5267 2748
rect 5267 2692 5271 2748
rect 5207 2688 5271 2692
rect 5287 2748 5351 2752
rect 5287 2692 5291 2748
rect 5291 2692 5347 2748
rect 5347 2692 5351 2748
rect 5287 2688 5351 2692
rect 5367 2748 5431 2752
rect 5367 2692 5371 2748
rect 5371 2692 5427 2748
rect 5427 2692 5431 2748
rect 5367 2688 5431 2692
rect 5447 2748 5511 2752
rect 5447 2692 5451 2748
rect 5451 2692 5507 2748
rect 5507 2692 5511 2748
rect 5447 2688 5511 2692
rect 6909 2748 6973 2752
rect 6909 2692 6913 2748
rect 6913 2692 6969 2748
rect 6969 2692 6973 2748
rect 6909 2688 6973 2692
rect 6989 2748 7053 2752
rect 6989 2692 6993 2748
rect 6993 2692 7049 2748
rect 7049 2692 7053 2748
rect 6989 2688 7053 2692
rect 7069 2748 7133 2752
rect 7069 2692 7073 2748
rect 7073 2692 7129 2748
rect 7129 2692 7133 2748
rect 7069 2688 7133 2692
rect 7149 2748 7213 2752
rect 7149 2692 7153 2748
rect 7153 2692 7209 2748
rect 7209 2692 7213 2748
rect 7149 2688 7213 2692
rect 2463 2204 2527 2208
rect 2463 2148 2467 2204
rect 2467 2148 2523 2204
rect 2523 2148 2527 2204
rect 2463 2144 2527 2148
rect 2543 2204 2607 2208
rect 2543 2148 2547 2204
rect 2547 2148 2603 2204
rect 2603 2148 2607 2204
rect 2543 2144 2607 2148
rect 2623 2204 2687 2208
rect 2623 2148 2627 2204
rect 2627 2148 2683 2204
rect 2683 2148 2687 2204
rect 2623 2144 2687 2148
rect 2703 2204 2767 2208
rect 2703 2148 2707 2204
rect 2707 2148 2763 2204
rect 2763 2148 2767 2204
rect 2703 2144 2767 2148
rect 4165 2204 4229 2208
rect 4165 2148 4169 2204
rect 4169 2148 4225 2204
rect 4225 2148 4229 2204
rect 4165 2144 4229 2148
rect 4245 2204 4309 2208
rect 4245 2148 4249 2204
rect 4249 2148 4305 2204
rect 4305 2148 4309 2204
rect 4245 2144 4309 2148
rect 4325 2204 4389 2208
rect 4325 2148 4329 2204
rect 4329 2148 4385 2204
rect 4385 2148 4389 2204
rect 4325 2144 4389 2148
rect 4405 2204 4469 2208
rect 4405 2148 4409 2204
rect 4409 2148 4465 2204
rect 4465 2148 4469 2204
rect 4405 2144 4469 2148
rect 5867 2204 5931 2208
rect 5867 2148 5871 2204
rect 5871 2148 5927 2204
rect 5927 2148 5931 2204
rect 5867 2144 5931 2148
rect 5947 2204 6011 2208
rect 5947 2148 5951 2204
rect 5951 2148 6007 2204
rect 6007 2148 6011 2204
rect 5947 2144 6011 2148
rect 6027 2204 6091 2208
rect 6027 2148 6031 2204
rect 6031 2148 6087 2204
rect 6087 2148 6091 2204
rect 6027 2144 6091 2148
rect 6107 2204 6171 2208
rect 6107 2148 6111 2204
rect 6111 2148 6167 2204
rect 6167 2148 6171 2204
rect 6107 2144 6171 2148
rect 7569 2204 7633 2208
rect 7569 2148 7573 2204
rect 7573 2148 7629 2204
rect 7629 2148 7633 2204
rect 7569 2144 7633 2148
rect 7649 2204 7713 2208
rect 7649 2148 7653 2204
rect 7653 2148 7709 2204
rect 7709 2148 7713 2204
rect 7649 2144 7713 2148
rect 7729 2204 7793 2208
rect 7729 2148 7733 2204
rect 7733 2148 7789 2204
rect 7789 2148 7793 2204
rect 7729 2144 7793 2148
rect 7809 2204 7873 2208
rect 7809 2148 7813 2204
rect 7813 2148 7869 2204
rect 7869 2148 7873 2204
rect 7809 2144 7873 2148
<< metal4 >>
rect 1795 8192 2115 8752
rect 1795 8128 1803 8192
rect 1867 8128 1883 8192
rect 1947 8128 1963 8192
rect 2027 8128 2043 8192
rect 2107 8128 2115 8192
rect 1795 8006 2115 8128
rect 1795 7770 1837 8006
rect 2073 7770 2115 8006
rect 1795 7104 2115 7770
rect 1795 7040 1803 7104
rect 1867 7040 1883 7104
rect 1947 7040 1963 7104
rect 2027 7040 2043 7104
rect 2107 7040 2115 7104
rect 1795 6374 2115 7040
rect 1795 6138 1837 6374
rect 2073 6138 2115 6374
rect 1795 6016 2115 6138
rect 1795 5952 1803 6016
rect 1867 5952 1883 6016
rect 1947 5952 1963 6016
rect 2027 5952 2043 6016
rect 2107 5952 2115 6016
rect 1795 4928 2115 5952
rect 1795 4864 1803 4928
rect 1867 4864 1883 4928
rect 1947 4864 1963 4928
rect 2027 4864 2043 4928
rect 2107 4864 2115 4928
rect 1795 4742 2115 4864
rect 1795 4506 1837 4742
rect 2073 4506 2115 4742
rect 1795 3840 2115 4506
rect 1795 3776 1803 3840
rect 1867 3776 1883 3840
rect 1947 3776 1963 3840
rect 2027 3776 2043 3840
rect 2107 3776 2115 3840
rect 1795 3110 2115 3776
rect 1795 2874 1837 3110
rect 2073 2874 2115 3110
rect 1795 2752 2115 2874
rect 1795 2688 1803 2752
rect 1867 2688 1883 2752
rect 1947 2688 1963 2752
rect 2027 2688 2043 2752
rect 2107 2688 2115 2752
rect 1795 2128 2115 2688
rect 2455 8736 2775 8752
rect 2455 8672 2463 8736
rect 2527 8672 2543 8736
rect 2607 8672 2623 8736
rect 2687 8672 2703 8736
rect 2767 8672 2775 8736
rect 2455 8666 2775 8672
rect 2455 8430 2497 8666
rect 2733 8430 2775 8666
rect 2455 7648 2775 8430
rect 2455 7584 2463 7648
rect 2527 7584 2543 7648
rect 2607 7584 2623 7648
rect 2687 7584 2703 7648
rect 2767 7584 2775 7648
rect 2455 7034 2775 7584
rect 2455 6798 2497 7034
rect 2733 6798 2775 7034
rect 2455 6560 2775 6798
rect 2455 6496 2463 6560
rect 2527 6496 2543 6560
rect 2607 6496 2623 6560
rect 2687 6496 2703 6560
rect 2767 6496 2775 6560
rect 2455 5472 2775 6496
rect 2455 5408 2463 5472
rect 2527 5408 2543 5472
rect 2607 5408 2623 5472
rect 2687 5408 2703 5472
rect 2767 5408 2775 5472
rect 2455 5402 2775 5408
rect 2455 5166 2497 5402
rect 2733 5166 2775 5402
rect 2455 4384 2775 5166
rect 2455 4320 2463 4384
rect 2527 4320 2543 4384
rect 2607 4320 2623 4384
rect 2687 4320 2703 4384
rect 2767 4320 2775 4384
rect 2455 3770 2775 4320
rect 2455 3534 2497 3770
rect 2733 3534 2775 3770
rect 2455 3296 2775 3534
rect 2455 3232 2463 3296
rect 2527 3232 2543 3296
rect 2607 3232 2623 3296
rect 2687 3232 2703 3296
rect 2767 3232 2775 3296
rect 2455 2208 2775 3232
rect 2455 2144 2463 2208
rect 2527 2144 2543 2208
rect 2607 2144 2623 2208
rect 2687 2144 2703 2208
rect 2767 2144 2775 2208
rect 2455 2128 2775 2144
rect 3497 8192 3817 8752
rect 3497 8128 3505 8192
rect 3569 8128 3585 8192
rect 3649 8128 3665 8192
rect 3729 8128 3745 8192
rect 3809 8128 3817 8192
rect 3497 8006 3817 8128
rect 3497 7770 3539 8006
rect 3775 7770 3817 8006
rect 3497 7104 3817 7770
rect 3497 7040 3505 7104
rect 3569 7040 3585 7104
rect 3649 7040 3665 7104
rect 3729 7040 3745 7104
rect 3809 7040 3817 7104
rect 3497 6374 3817 7040
rect 3497 6138 3539 6374
rect 3775 6138 3817 6374
rect 3497 6016 3817 6138
rect 3497 5952 3505 6016
rect 3569 5952 3585 6016
rect 3649 5952 3665 6016
rect 3729 5952 3745 6016
rect 3809 5952 3817 6016
rect 3497 4928 3817 5952
rect 3497 4864 3505 4928
rect 3569 4864 3585 4928
rect 3649 4864 3665 4928
rect 3729 4864 3745 4928
rect 3809 4864 3817 4928
rect 3497 4742 3817 4864
rect 3497 4506 3539 4742
rect 3775 4506 3817 4742
rect 3497 3840 3817 4506
rect 3497 3776 3505 3840
rect 3569 3776 3585 3840
rect 3649 3776 3665 3840
rect 3729 3776 3745 3840
rect 3809 3776 3817 3840
rect 3497 3110 3817 3776
rect 3497 2874 3539 3110
rect 3775 2874 3817 3110
rect 3497 2752 3817 2874
rect 3497 2688 3505 2752
rect 3569 2688 3585 2752
rect 3649 2688 3665 2752
rect 3729 2688 3745 2752
rect 3809 2688 3817 2752
rect 3497 2128 3817 2688
rect 4157 8736 4477 8752
rect 4157 8672 4165 8736
rect 4229 8672 4245 8736
rect 4309 8672 4325 8736
rect 4389 8672 4405 8736
rect 4469 8672 4477 8736
rect 4157 8666 4477 8672
rect 4157 8430 4199 8666
rect 4435 8430 4477 8666
rect 4157 7648 4477 8430
rect 4157 7584 4165 7648
rect 4229 7584 4245 7648
rect 4309 7584 4325 7648
rect 4389 7584 4405 7648
rect 4469 7584 4477 7648
rect 4157 7034 4477 7584
rect 4157 6798 4199 7034
rect 4435 6798 4477 7034
rect 4157 6560 4477 6798
rect 4157 6496 4165 6560
rect 4229 6496 4245 6560
rect 4309 6496 4325 6560
rect 4389 6496 4405 6560
rect 4469 6496 4477 6560
rect 4157 5472 4477 6496
rect 4157 5408 4165 5472
rect 4229 5408 4245 5472
rect 4309 5408 4325 5472
rect 4389 5408 4405 5472
rect 4469 5408 4477 5472
rect 4157 5402 4477 5408
rect 4157 5166 4199 5402
rect 4435 5166 4477 5402
rect 4157 4384 4477 5166
rect 4157 4320 4165 4384
rect 4229 4320 4245 4384
rect 4309 4320 4325 4384
rect 4389 4320 4405 4384
rect 4469 4320 4477 4384
rect 4157 3770 4477 4320
rect 4157 3534 4199 3770
rect 4435 3534 4477 3770
rect 4157 3296 4477 3534
rect 4157 3232 4165 3296
rect 4229 3232 4245 3296
rect 4309 3232 4325 3296
rect 4389 3232 4405 3296
rect 4469 3232 4477 3296
rect 4157 2208 4477 3232
rect 4157 2144 4165 2208
rect 4229 2144 4245 2208
rect 4309 2144 4325 2208
rect 4389 2144 4405 2208
rect 4469 2144 4477 2208
rect 4157 2128 4477 2144
rect 5199 8192 5519 8752
rect 5199 8128 5207 8192
rect 5271 8128 5287 8192
rect 5351 8128 5367 8192
rect 5431 8128 5447 8192
rect 5511 8128 5519 8192
rect 5199 8006 5519 8128
rect 5199 7770 5241 8006
rect 5477 7770 5519 8006
rect 5199 7104 5519 7770
rect 5199 7040 5207 7104
rect 5271 7040 5287 7104
rect 5351 7040 5367 7104
rect 5431 7040 5447 7104
rect 5511 7040 5519 7104
rect 5199 6374 5519 7040
rect 5199 6138 5241 6374
rect 5477 6138 5519 6374
rect 5199 6016 5519 6138
rect 5199 5952 5207 6016
rect 5271 5952 5287 6016
rect 5351 5952 5367 6016
rect 5431 5952 5447 6016
rect 5511 5952 5519 6016
rect 5199 4928 5519 5952
rect 5199 4864 5207 4928
rect 5271 4864 5287 4928
rect 5351 4864 5367 4928
rect 5431 4864 5447 4928
rect 5511 4864 5519 4928
rect 5199 4742 5519 4864
rect 5199 4506 5241 4742
rect 5477 4506 5519 4742
rect 5199 3840 5519 4506
rect 5199 3776 5207 3840
rect 5271 3776 5287 3840
rect 5351 3776 5367 3840
rect 5431 3776 5447 3840
rect 5511 3776 5519 3840
rect 5199 3110 5519 3776
rect 5199 2874 5241 3110
rect 5477 2874 5519 3110
rect 5199 2752 5519 2874
rect 5199 2688 5207 2752
rect 5271 2688 5287 2752
rect 5351 2688 5367 2752
rect 5431 2688 5447 2752
rect 5511 2688 5519 2752
rect 5199 2128 5519 2688
rect 5859 8736 6179 8752
rect 5859 8672 5867 8736
rect 5931 8672 5947 8736
rect 6011 8672 6027 8736
rect 6091 8672 6107 8736
rect 6171 8672 6179 8736
rect 5859 8666 6179 8672
rect 5859 8430 5901 8666
rect 6137 8430 6179 8666
rect 5859 7648 6179 8430
rect 5859 7584 5867 7648
rect 5931 7584 5947 7648
rect 6011 7584 6027 7648
rect 6091 7584 6107 7648
rect 6171 7584 6179 7648
rect 5859 7034 6179 7584
rect 5859 6798 5901 7034
rect 6137 6798 6179 7034
rect 5859 6560 6179 6798
rect 5859 6496 5867 6560
rect 5931 6496 5947 6560
rect 6011 6496 6027 6560
rect 6091 6496 6107 6560
rect 6171 6496 6179 6560
rect 5859 5472 6179 6496
rect 5859 5408 5867 5472
rect 5931 5408 5947 5472
rect 6011 5408 6027 5472
rect 6091 5408 6107 5472
rect 6171 5408 6179 5472
rect 5859 5402 6179 5408
rect 5859 5166 5901 5402
rect 6137 5166 6179 5402
rect 5859 4384 6179 5166
rect 5859 4320 5867 4384
rect 5931 4320 5947 4384
rect 6011 4320 6027 4384
rect 6091 4320 6107 4384
rect 6171 4320 6179 4384
rect 5859 3770 6179 4320
rect 5859 3534 5901 3770
rect 6137 3534 6179 3770
rect 5859 3296 6179 3534
rect 5859 3232 5867 3296
rect 5931 3232 5947 3296
rect 6011 3232 6027 3296
rect 6091 3232 6107 3296
rect 6171 3232 6179 3296
rect 5859 2208 6179 3232
rect 5859 2144 5867 2208
rect 5931 2144 5947 2208
rect 6011 2144 6027 2208
rect 6091 2144 6107 2208
rect 6171 2144 6179 2208
rect 5859 2128 6179 2144
rect 6901 8192 7221 8752
rect 6901 8128 6909 8192
rect 6973 8128 6989 8192
rect 7053 8128 7069 8192
rect 7133 8128 7149 8192
rect 7213 8128 7221 8192
rect 6901 8006 7221 8128
rect 6901 7770 6943 8006
rect 7179 7770 7221 8006
rect 6901 7104 7221 7770
rect 6901 7040 6909 7104
rect 6973 7040 6989 7104
rect 7053 7040 7069 7104
rect 7133 7040 7149 7104
rect 7213 7040 7221 7104
rect 6901 6374 7221 7040
rect 6901 6138 6943 6374
rect 7179 6138 7221 6374
rect 6901 6016 7221 6138
rect 6901 5952 6909 6016
rect 6973 5952 6989 6016
rect 7053 5952 7069 6016
rect 7133 5952 7149 6016
rect 7213 5952 7221 6016
rect 6901 4928 7221 5952
rect 6901 4864 6909 4928
rect 6973 4864 6989 4928
rect 7053 4864 7069 4928
rect 7133 4864 7149 4928
rect 7213 4864 7221 4928
rect 6901 4742 7221 4864
rect 6901 4506 6943 4742
rect 7179 4506 7221 4742
rect 6901 3840 7221 4506
rect 6901 3776 6909 3840
rect 6973 3776 6989 3840
rect 7053 3776 7069 3840
rect 7133 3776 7149 3840
rect 7213 3776 7221 3840
rect 6901 3110 7221 3776
rect 6901 2874 6943 3110
rect 7179 2874 7221 3110
rect 6901 2752 7221 2874
rect 6901 2688 6909 2752
rect 6973 2688 6989 2752
rect 7053 2688 7069 2752
rect 7133 2688 7149 2752
rect 7213 2688 7221 2752
rect 6901 2128 7221 2688
rect 7561 8736 7881 8752
rect 7561 8672 7569 8736
rect 7633 8672 7649 8736
rect 7713 8672 7729 8736
rect 7793 8672 7809 8736
rect 7873 8672 7881 8736
rect 7561 8666 7881 8672
rect 7561 8430 7603 8666
rect 7839 8430 7881 8666
rect 7561 7648 7881 8430
rect 7561 7584 7569 7648
rect 7633 7584 7649 7648
rect 7713 7584 7729 7648
rect 7793 7584 7809 7648
rect 7873 7584 7881 7648
rect 7561 7034 7881 7584
rect 7561 6798 7603 7034
rect 7839 6798 7881 7034
rect 7561 6560 7881 6798
rect 7561 6496 7569 6560
rect 7633 6496 7649 6560
rect 7713 6496 7729 6560
rect 7793 6496 7809 6560
rect 7873 6496 7881 6560
rect 7561 5472 7881 6496
rect 7561 5408 7569 5472
rect 7633 5408 7649 5472
rect 7713 5408 7729 5472
rect 7793 5408 7809 5472
rect 7873 5408 7881 5472
rect 7561 5402 7881 5408
rect 7561 5166 7603 5402
rect 7839 5166 7881 5402
rect 7561 4384 7881 5166
rect 7561 4320 7569 4384
rect 7633 4320 7649 4384
rect 7713 4320 7729 4384
rect 7793 4320 7809 4384
rect 7873 4320 7881 4384
rect 7561 3770 7881 4320
rect 7561 3534 7603 3770
rect 7839 3534 7881 3770
rect 7561 3296 7881 3534
rect 7561 3232 7569 3296
rect 7633 3232 7649 3296
rect 7713 3232 7729 3296
rect 7793 3232 7809 3296
rect 7873 3232 7881 3296
rect 7561 2208 7881 3232
rect 7561 2144 7569 2208
rect 7633 2144 7649 2208
rect 7713 2144 7729 2208
rect 7793 2144 7809 2208
rect 7873 2144 7881 2208
rect 7561 2128 7881 2144
<< via4 >>
rect 1837 7770 2073 8006
rect 1837 6138 2073 6374
rect 1837 4506 2073 4742
rect 1837 2874 2073 3110
rect 2497 8430 2733 8666
rect 2497 6798 2733 7034
rect 2497 5166 2733 5402
rect 2497 3534 2733 3770
rect 3539 7770 3775 8006
rect 3539 6138 3775 6374
rect 3539 4506 3775 4742
rect 3539 2874 3775 3110
rect 4199 8430 4435 8666
rect 4199 6798 4435 7034
rect 4199 5166 4435 5402
rect 4199 3534 4435 3770
rect 5241 7770 5477 8006
rect 5241 6138 5477 6374
rect 5241 4506 5477 4742
rect 5241 2874 5477 3110
rect 5901 8430 6137 8666
rect 5901 6798 6137 7034
rect 5901 5166 6137 5402
rect 5901 3534 6137 3770
rect 6943 7770 7179 8006
rect 6943 6138 7179 6374
rect 6943 4506 7179 4742
rect 6943 2874 7179 3110
rect 7603 8430 7839 8666
rect 7603 6798 7839 7034
rect 7603 5166 7839 5402
rect 7603 3534 7839 3770
<< metal5 >>
rect 1056 8666 7960 8708
rect 1056 8430 2497 8666
rect 2733 8430 4199 8666
rect 4435 8430 5901 8666
rect 6137 8430 7603 8666
rect 7839 8430 7960 8666
rect 1056 8388 7960 8430
rect 1056 8006 7960 8048
rect 1056 7770 1837 8006
rect 2073 7770 3539 8006
rect 3775 7770 5241 8006
rect 5477 7770 6943 8006
rect 7179 7770 7960 8006
rect 1056 7728 7960 7770
rect 1056 7034 7960 7076
rect 1056 6798 2497 7034
rect 2733 6798 4199 7034
rect 4435 6798 5901 7034
rect 6137 6798 7603 7034
rect 7839 6798 7960 7034
rect 1056 6756 7960 6798
rect 1056 6374 7960 6416
rect 1056 6138 1837 6374
rect 2073 6138 3539 6374
rect 3775 6138 5241 6374
rect 5477 6138 6943 6374
rect 7179 6138 7960 6374
rect 1056 6096 7960 6138
rect 1056 5402 7960 5444
rect 1056 5166 2497 5402
rect 2733 5166 4199 5402
rect 4435 5166 5901 5402
rect 6137 5166 7603 5402
rect 7839 5166 7960 5402
rect 1056 5124 7960 5166
rect 1056 4742 7960 4784
rect 1056 4506 1837 4742
rect 2073 4506 3539 4742
rect 3775 4506 5241 4742
rect 5477 4506 6943 4742
rect 7179 4506 7960 4742
rect 1056 4464 7960 4506
rect 1056 3770 7960 3812
rect 1056 3534 2497 3770
rect 2733 3534 4199 3770
rect 4435 3534 5901 3770
rect 6137 3534 7603 3770
rect 7839 3534 7960 3770
rect 1056 3492 7960 3534
rect 1056 3110 7960 3152
rect 1056 2874 1837 3110
rect 2073 2874 3539 3110
rect 3775 2874 5241 3110
rect 5477 2874 6943 3110
rect 7179 2874 7960 3110
rect 1056 2832 7960 2874
use sky130_fd_sc_hd__buf_2  _34_ ~/Openlane/install/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1698771642
transform 1 0 4508 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _35_
timestamp 1698771642
transform 1 0 4324 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__nor3b_1  _36_ ~/Openlane/install/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1698771642
transform 1 0 3772 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_2  _37_ ~/Openlane/install/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1698771642
transform 1 0 2668 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__buf_2  _38_
timestamp 1698771642
transform -1 0 2668 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _39_ ~/Openlane/install/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1698771642
transform 1 0 1472 0 -1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _40_ ~/Openlane/install/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1698771642
transform 1 0 2208 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__o31a_1  _41_ ~/Openlane/install/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1698771642
transform -1 0 3312 0 1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__nor3b_1  _42_
timestamp 1698771642
transform 1 0 6900 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  _43_ ~/Openlane/install/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1698771642
transform 1 0 5520 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _44_
timestamp 1698771642
transform 1 0 4876 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__o31a_1  _45_
timestamp 1698771642
transform 1 0 4600 0 -1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__nor3b_1  _46_
timestamp 1698771642
transform 1 0 6348 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  _47_
timestamp 1698771642
transform -1 0 5888 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _48_
timestamp 1698771642
transform 1 0 4876 0 1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__o31a_1  _49_
timestamp 1698771642
transform -1 0 5888 0 -1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__nor3b_1  _50_
timestamp 1698771642
transform -1 0 4048 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  _51_
timestamp 1698771642
transform 1 0 4140 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _52_
timestamp 1698771642
transform 1 0 3772 0 1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__o31a_1  _53_
timestamp 1698771642
transform 1 0 3772 0 -1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__nor3b_1  _54_
timestamp 1698771642
transform 1 0 3404 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  _55_
timestamp 1698771642
transform 1 0 3128 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _56_
timestamp 1698771642
transform 1 0 2668 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__o31a_1  _57_
timestamp 1698771642
transform 1 0 2668 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__nor3b_1  _58_
timestamp 1698771642
transform 1 0 4140 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  _59_
timestamp 1698771642
transform 1 0 3956 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _60_
timestamp 1698771642
transform 1 0 4048 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__o31a_1  _61_
timestamp 1698771642
transform 1 0 3772 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__nor3b_1  _62_
timestamp 1698771642
transform 1 0 4968 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  _63_
timestamp 1698771642
transform -1 0 5336 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _64_
timestamp 1698771642
transform 1 0 4416 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__o31a_1  _65_
timestamp 1698771642
transform -1 0 5520 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _66_ ~/Openlane/install/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1698771642
transform -1 0 5244 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__o32a_1  _67_ ~/Openlane/install/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1698771642
transform 1 0 6348 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dfrtp_1  _68_ ~/Openlane/install/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1698771642
transform 1 0 1748 0 1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _69_
timestamp 1698771642
transform 1 0 5336 0 1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _70_
timestamp 1698771642
transform 1 0 5336 0 1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _71_
timestamp 1698771642
transform 1 0 1932 0 -1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _72_
timestamp 1698771642
transform -1 0 3404 0 1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _73_
timestamp 1698771642
transform 1 0 2300 0 -1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _74_
timestamp 1698771642
transform 1 0 5244 0 1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _75_
timestamp 1698771642
transform 1 0 5520 0 1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_1  _76_ ~/Openlane/install/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1698771642
transform 1 0 7360 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_clk ~/Openlane/install/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1698771642
transform 1 0 3772 0 1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_0__f_clk
timestamp 1698771642
transform -1 0 4600 0 -1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_1__f_clk
timestamp 1698771642
transform -1 0 3680 0 -1 8704
box -38 -48 1878 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_3 ~/Openlane/install/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1698771642
transform 1 0 1380 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_15
timestamp 1698771642
transform 1 0 2484 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_27 ~/Openlane/install/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1698771642
transform 1 0 3588 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_34
timestamp 1698771642
transform 1 0 4232 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_46 ~/Openlane/install/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1698771642
transform 1 0 5336 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_54 ~/Openlane/install/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1698771642
transform 1 0 6072 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_0_57 ~/Openlane/install/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1698771642
transform 1 0 6348 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_69
timestamp 1698771642
transform 1 0 7452 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_13 ~/Openlane/install/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1698771642
transform 1 0 2300 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_17
timestamp 1698771642
transform 1 0 2668 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1_38
timestamp 1698771642
transform 1 0 4600 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_46
timestamp 1698771642
transform 1 0 5336 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_54
timestamp 1698771642
transform 1 0 6072 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_65
timestamp 1698771642
transform 1 0 7084 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2_3
timestamp 1698771642
transform 1 0 1380 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_27
timestamp 1698771642
transform 1 0 3588 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2_29
timestamp 1698771642
transform 1 0 3772 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_39
timestamp 1698771642
transform 1 0 4692 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_66
timestamp 1698771642
transform 1 0 7176 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_3
timestamp 1698771642
transform 1 0 1380 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_36
timestamp 1698771642
transform 1 0 4416 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_52
timestamp 1698771642
transform 1 0 5888 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_69
timestamp 1698771642
transform 1 0 7452 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_4_3
timestamp 1698771642
transform 1 0 1380 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_11
timestamp 1698771642
transform 1 0 2116 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_4_24
timestamp 1698771642
transform 1 0 3312 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_39
timestamp 1698771642
transform 1 0 4692 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_66
timestamp 1698771642
transform 1 0 7176 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_6
timestamp 1698771642
transform 1 0 1656 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_5_18
timestamp 1698771642
transform 1 0 2760 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_5_37
timestamp 1698771642
transform 1 0 4508 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_45
timestamp 1698771642
transform 1 0 5244 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_52
timestamp 1698771642
transform 1 0 5888 0 -1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_57
timestamp 1698771642
transform 1 0 6348 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_69
timestamp 1698771642
transform 1 0 7452 0 -1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_3
timestamp 1698771642
transform 1 0 1380 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_15
timestamp 1698771642
transform 1 0 2484 0 1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_49
timestamp 1698771642
transform 1 0 5612 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_6_61
timestamp 1698771642
transform 1 0 6716 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_7
timestamp 1698771642
transform 1 0 1748 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_24
timestamp 1698771642
transform 1 0 3312 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_7_37 ~/Openlane/install/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1698771642
transform 1 0 4508 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_7_46
timestamp 1698771642
transform 1 0 5336 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_54
timestamp 1698771642
transform 1 0 6072 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_65
timestamp 1698771642
transform 1 0 7084 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_3
timestamp 1698771642
transform 1 0 1380 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_8_25
timestamp 1698771642
transform 1 0 3404 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_9_3
timestamp 1698771642
transform 1 0 1380 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_11
timestamp 1698771642
transform 1 0 2116 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_9_39
timestamp 1698771642
transform 1 0 4692 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_10_9
timestamp 1698771642
transform 1 0 1932 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_22
timestamp 1698771642
transform 1 0 3128 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_10_29
timestamp 1698771642
transform 1 0 3772 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_65
timestamp 1698771642
transform 1 0 7084 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_3
timestamp 1698771642
transform 1 0 1380 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_29
timestamp 1698771642
transform 1 0 3772 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_41
timestamp 1698771642
transform 1 0 4876 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_11_53
timestamp 1698771642
transform 1 0 5980 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold1 ~/Openlane/install/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1698771642
transform -1 0 7636 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold2
timestamp 1698771642
transform -1 0 6256 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold3
timestamp 1698771642
transform -1 0 7084 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold4
timestamp 1698771642
transform -1 0 7084 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  input1
timestamp 1698771642
transform 1 0 1472 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  input2 ~/Openlane/install/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1698771642
transform 1 0 1380 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  input3 ~/Openlane/install/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1698771642
transform 1 0 1380 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input4
timestamp 1698771642
transform -1 0 1656 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input5 ~/Openlane/install/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1698771642
transform 1 0 1380 0 -1 3264
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_4  output6
timestamp 1698771642
transform 1 0 6900 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output7
timestamp 1698771642
transform 1 0 7268 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output8
timestamp 1698771642
transform 1 0 7268 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output9
timestamp 1698771642
transform 1 0 7268 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output10
timestamp 1698771642
transform 1 0 7084 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output11
timestamp 1698771642
transform 1 0 7268 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output12
timestamp 1698771642
transform 1 0 7268 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output13
timestamp 1698771642
transform 1 0 7084 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output14
timestamp 1698771642
transform -1 0 6900 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Left_12
timestamp 1698771642
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Right_0
timestamp 1698771642
transform -1 0 7912 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Left_13
timestamp 1698771642
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Right_1
timestamp 1698771642
transform -1 0 7912 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Left_14
timestamp 1698771642
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Right_2
timestamp 1698771642
transform -1 0 7912 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Left_15
timestamp 1698771642
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Right_3
timestamp 1698771642
transform -1 0 7912 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Left_16
timestamp 1698771642
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Right_4
timestamp 1698771642
transform -1 0 7912 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Left_17
timestamp 1698771642
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Right_5
timestamp 1698771642
transform -1 0 7912 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Left_18
timestamp 1698771642
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Right_6
timestamp 1698771642
transform -1 0 7912 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Left_19
timestamp 1698771642
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Right_7
timestamp 1698771642
transform -1 0 7912 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Left_20
timestamp 1698771642
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Right_8
timestamp 1698771642
transform -1 0 7912 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Left_21
timestamp 1698771642
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Right_9
timestamp 1698771642
transform -1 0 7912 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_Left_22
timestamp 1698771642
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_Right_10
timestamp 1698771642
transform -1 0 7912 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_Left_23
timestamp 1698771642
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_Right_11
timestamp 1698771642
transform -1 0 7912 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_24 ~/Openlane/install/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1698771642
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_25
timestamp 1698771642
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_26
timestamp 1698771642
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_27
timestamp 1698771642
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_28
timestamp 1698771642
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_29
timestamp 1698771642
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_30
timestamp 1698771642
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_31
timestamp 1698771642
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_32
timestamp 1698771642
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_33
timestamp 1698771642
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_34
timestamp 1698771642
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_35
timestamp 1698771642
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_36
timestamp 1698771642
transform 1 0 3680 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_37
timestamp 1698771642
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
<< labels >>
flabel metal4 s 2455 2128 2775 8752 0 FreeSans 1920 90 0 0 GND
port 0 nsew ground bidirectional
flabel metal4 s 4157 2128 4477 8752 0 FreeSans 1920 90 0 0 GND
port 0 nsew ground bidirectional
flabel metal4 s 5859 2128 6179 8752 0 FreeSans 1920 90 0 0 GND
port 0 nsew ground bidirectional
flabel metal4 s 7561 2128 7881 8752 0 FreeSans 1920 90 0 0 GND
port 0 nsew ground bidirectional
flabel metal5 s 1056 3492 7960 3812 0 FreeSans 2560 0 0 0 GND
port 0 nsew ground bidirectional
flabel metal5 s 1056 5124 7960 5444 0 FreeSans 2560 0 0 0 GND
port 0 nsew ground bidirectional
flabel metal5 s 1056 6756 7960 7076 0 FreeSans 2560 0 0 0 GND
port 0 nsew ground bidirectional
flabel metal5 s 1056 8388 7960 8708 0 FreeSans 2560 0 0 0 GND
port 0 nsew ground bidirectional
flabel metal4 s 1795 2128 2115 8752 0 FreeSans 1920 90 0 0 VDD
port 1 nsew power bidirectional
flabel metal4 s 3497 2128 3817 8752 0 FreeSans 1920 90 0 0 VDD
port 1 nsew power bidirectional
flabel metal4 s 5199 2128 5519 8752 0 FreeSans 1920 90 0 0 VDD
port 1 nsew power bidirectional
flabel metal4 s 6901 2128 7221 8752 0 FreeSans 1920 90 0 0 VDD
port 1 nsew power bidirectional
flabel metal5 s 1056 2832 7960 3152 0 FreeSans 2560 0 0 0 VDD
port 1 nsew power bidirectional
flabel metal5 s 1056 4464 7960 4784 0 FreeSans 2560 0 0 0 VDD
port 1 nsew power bidirectional
flabel metal5 s 1056 6096 7960 6416 0 FreeSans 2560 0 0 0 VDD
port 1 nsew power bidirectional
flabel metal5 s 1056 7728 7960 8048 0 FreeSans 2560 0 0 0 VDD
port 1 nsew power bidirectional
flabel metal3 s 8226 1096 9026 1216 0 FreeSans 480 0 0 0 data_out[0]
port 3 nsew signal tristate
flabel metal3 s 8226 2184 9026 2304 0 FreeSans 480 0 0 0 data_out[1]
port 4 nsew signal tristate
flabel metal3 s 8226 3272 9026 3392 0 FreeSans 480 0 0 0 data_out[2]
port 5 nsew signal tristate
flabel metal3 s 8226 4360 9026 4480 0 FreeSans 480 0 0 0 data_out[3]
port 6 nsew signal tristate
flabel metal3 s 8226 5448 9026 5568 0 FreeSans 480 0 0 0 data_out[4]
port 7 nsew signal tristate
flabel metal3 s 8226 6536 9026 6656 0 FreeSans 480 0 0 0 data_out[5]
port 8 nsew signal tristate
flabel metal3 s 8226 7624 9026 7744 0 FreeSans 480 0 0 0 data_out[6]
port 9 nsew signal tristate
flabel metal3 s 8226 8712 9026 8832 0 FreeSans 480 0 0 0 data_out[7]
port 10 nsew signal tristate
flabel metal3 s 8226 9800 9026 9920 0 FreeSans 480 0 0 0 scan_out
port 15 nsew signal tristate
rlabel metal1 4508 8704 4508 8704 0 GND
rlabel metal1 4508 8160 4508 8160 0 VDD
rlabel metal1 2070 3400 2070 3400 0 _00_
rlabel metal1 5152 4250 5152 4250 0 _01_
rlabel metal1 5704 3570 5704 3570 0 _02_
rlabel metal1 3036 4046 3036 4046 0 _03_
rlabel metal2 3082 6562 3082 6562 0 _04_
rlabel metal1 3588 6698 3588 6698 0 _05_
rlabel metal1 5612 6698 5612 6698 0 _06_
rlabel metal2 6394 6868 6394 6868 0 _07_
rlabel metal1 6808 4046 6808 4046 0 _08_
rlabel metal2 6578 3502 6578 3502 0 _09_
rlabel metal1 3450 4590 3450 4590 0 _10_
rlabel metal1 2898 6324 2898 6324 0 _11_
rlabel metal2 2346 5372 2346 5372 0 _12_
rlabel metal2 2990 4318 2990 4318 0 _13_
rlabel metal1 2622 4522 2622 4522 0 _14_
rlabel metal1 4968 4114 4968 4114 0 _15_
rlabel metal1 5244 3162 5244 3162 0 _16_
rlabel metal1 5198 4114 5198 4114 0 _17_
rlabel metal1 5980 3978 5980 3978 0 _18_
rlabel metal1 5520 4114 5520 4114 0 _19_
rlabel metal1 5336 3706 5336 3706 0 _20_
rlabel metal1 4048 3978 4048 3978 0 _21_
rlabel metal2 4186 3842 4186 3842 0 _22_
rlabel metal1 4416 2618 4416 2618 0 _23_
rlabel metal1 3220 6222 3220 6222 0 _24_
rlabel metal1 3128 5882 3128 5882 0 _25_
rlabel metal1 3128 5542 3128 5542 0 _26_
rlabel metal1 4140 6834 4140 6834 0 _27_
rlabel metal1 4048 6426 4048 6426 0 _28_
rlabel metal1 4508 5338 4508 5338 0 _29_
rlabel metal1 5106 6902 5106 6902 0 _30_
rlabel metal1 5244 6426 5244 6426 0 _31_
rlabel metal1 4922 6766 4922 6766 0 _32_
rlabel metal1 6992 6290 6992 6290 0 _33_
rlabel metal2 5106 7174 5106 7174 0 clknet_0_clk
rlabel metal1 5336 3570 5336 3570 0 clknet_1_0__leaf_clk
rlabel metal2 2346 7820 2346 7820 0 clknet_1_1__leaf_clk
rlabel metal1 6992 2278 6992 2278 0 data_out[0]
rlabel metal3 8196 2244 8196 2244 0 data_out[1]
rlabel metal1 7774 3366 7774 3366 0 data_out[2]
rlabel metal1 7774 4454 7774 4454 0 data_out[3]
rlabel metal1 7774 5542 7774 5542 0 data_out[4]
rlabel metal1 7774 6426 7774 6426 0 data_out[5]
rlabel metal1 7774 7718 7774 7718 0 data_out[6]
rlabel metal1 7728 7514 7728 7514 0 data_out[7]
rlabel metal2 2898 8092 2898 8092 0 net1
rlabel metal1 4232 6290 4232 6290 0 net10
rlabel metal1 5796 6290 5796 6290 0 net11
rlabel metal2 6946 7378 6946 7378 0 net12
rlabel metal1 6302 7378 6302 7378 0 net13
rlabel metal2 7406 7548 7406 7548 0 net14
rlabel metal1 6854 6324 6854 6324 0 net15
rlabel metal1 5740 6970 5740 6970 0 net16
rlabel metal1 6026 3162 6026 3162 0 net17
rlabel metal1 4462 6800 4462 6800 0 net18
rlabel metal1 1787 6766 1787 6766 0 net2
rlabel metal1 2162 6290 2162 6290 0 net3
rlabel metal1 1656 4114 1656 4114 0 net4
rlabel metal2 4554 3230 4554 3230 0 net5
rlabel metal1 2254 4658 2254 4658 0 net6
rlabel metal1 7268 4454 7268 4454 0 net7
rlabel metal1 5750 3366 5750 3366 0 net8
rlabel metal1 3542 3978 3542 3978 0 net9
rlabel metal1 1242 7854 1242 7854 0 reset
rlabel metal2 6670 9231 6670 9231 0 scan_out
<< properties >>
string FIXED_BBOX 0 0 9026 11170
<< end >>
