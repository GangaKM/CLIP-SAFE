magic
tech sky130A
magscale 1 2
timestamp 1698476459
<< error_s >>
rect 130 1084 192 1336
rect 222 1084 288 1336
rect 318 1084 384 1336
rect 414 1084 480 1336
rect 510 1084 576 1336
rect 606 1084 672 1336
rect 702 1084 768 1336
rect 798 1084 864 1336
rect 894 1084 960 1336
rect 990 1084 1056 1336
rect 1086 1084 1152 1336
rect 1182 1084 1248 1336
rect 1278 1084 1344 1336
rect 1374 1084 1440 1336
rect 1470 1084 1536 1336
rect 1566 1084 1632 1336
rect 1662 1084 1728 1336
rect 1758 1084 1824 1336
rect 1854 1084 1920 1336
rect 1950 1084 2016 1336
rect 2046 1084 2112 1336
rect 2142 1084 2208 1336
rect 2238 1084 2304 1336
rect 2334 1084 2400 1336
rect 2430 1084 2496 1336
rect 2526 1084 2579 1336
rect 130 622 192 706
rect 222 622 288 706
rect 318 622 384 706
rect 414 622 480 706
rect 510 622 576 706
rect 606 622 672 706
rect 702 622 768 706
rect 798 622 864 706
rect 894 622 960 706
rect 990 622 1056 706
rect 1086 622 1152 706
rect 1182 622 1248 706
rect 1278 622 1344 706
rect 1374 622 1440 706
rect 1470 622 1536 706
rect 1566 622 1632 706
rect 1662 622 1728 706
rect 1758 622 1824 706
rect 1854 622 1920 706
rect 1950 622 2016 706
rect 2046 622 2112 706
rect 2142 622 2208 706
rect 2238 622 2304 706
rect 2334 622 2400 706
rect 2430 622 2496 706
rect 2526 622 2585 706
<< nwell >>
rect 5326 1434 5686 1444
rect 5326 1416 5752 1434
rect 5388 1372 5752 1416
<< poly >>
rect -88 846 226 860
rect -88 790 -64 846
rect 198 790 226 846
rect -88 772 226 790
<< polycont >>
rect -64 790 198 846
<< locali >>
rect -88 846 226 860
rect -88 790 -64 846
rect 198 790 226 846
rect -88 772 226 790
<< viali >>
rect -64 790 198 846
<< metal1 >>
rect 3956 2014 4964 2020
rect 4 1968 4964 2014
rect 4 1476 120 1968
rect 4836 1476 4964 1968
rect 4 1444 4964 1476
rect 7086 880 7162 914
rect 5444 870 5472 874
rect 6166 870 6294 874
rect -88 846 226 860
rect -88 790 -64 846
rect 198 790 226 846
rect 5444 838 6294 870
rect 5446 820 6294 838
rect -88 772 226 790
rect 110 526 5386 534
rect 110 452 136 526
rect 5360 452 5386 526
rect 110 444 5386 452
<< via1 >>
rect 120 1476 4836 1968
rect -64 790 198 846
rect 136 452 5360 526
<< metal2 >>
rect 3956 2014 4964 2020
rect 4 1968 4964 2014
rect 4 1476 120 1968
rect 4836 1476 4964 1968
rect 4 1444 4964 1476
rect -84 918 5640 958
rect -88 846 226 860
rect -88 790 -64 846
rect 198 790 226 846
rect -88 772 226 790
rect 110 526 5386 534
rect 110 452 136 526
rect 5360 452 5386 526
rect 110 444 5386 452
<< via2 >>
rect 120 1504 4836 1940
rect -64 790 198 846
rect 136 452 5360 526
<< metal3 >>
rect 3956 2014 4964 2020
rect 4 1968 4964 2014
rect 4 1476 120 1968
rect 4836 1476 4964 1968
rect 4 1444 4964 1476
rect -116 846 226 860
rect -116 790 -64 846
rect 198 790 226 846
rect -116 772 226 790
rect -116 770 -54 772
rect 110 528 5386 534
rect 110 452 136 528
rect 474 526 5386 528
rect 5360 452 5386 526
rect 110 444 5386 452
<< via3 >>
rect 120 1940 4836 1968
rect 120 1504 4836 1940
rect 120 1476 4836 1504
rect 136 526 474 528
rect 136 452 5360 526
<< metal4 >>
rect 3956 2016 5700 2020
rect 3956 2014 6118 2016
rect 4 1968 7470 2014
rect 4 1476 120 1968
rect 4836 1476 7470 1968
rect 4 1444 7470 1476
rect 5110 1440 7470 1444
rect 5620 1434 7470 1440
rect 8 528 5504 540
rect 8 452 136 528
rect 474 526 5504 528
rect 5360 452 5504 526
rect 8 434 5504 452
rect 8 90 136 434
rect 4804 90 5504 434
rect 8 -2 5504 90
<< via4 >>
rect 136 90 4804 434
<< metal5 >>
rect -8 540 5504 544
rect -8 434 7448 540
rect -8 90 136 434
rect 4804 90 7448 434
rect -8 -30 7448 90
use and_gate  and_gate_0 ~/Desktop/charge_pumps2/layout_files
timestamp 1698389451
transform 1 0 5762 0 1 690
box -684 -688 1688 1316
use buffer  buffer_0 ~/Desktop/charge_pumps2/layout_files
timestamp 1698060067
transform 1 0 1330 0 1 -776
box -1330 776 4190 2342
<< labels >>
rlabel metal2 82 938 82 938 1 in1
port 1 n
rlabel metal3 -106 818 -106 818 1 clk
port 2 n
rlabel via4 4616 242 4616 242 1 gnd
port 3 n
rlabel metal4 5346 1798 5346 1798 1 vdd
port 4 n
rlabel metal1 7102 888 7102 888 1 out
port 5 n
<< end >>
