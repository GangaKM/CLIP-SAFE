magic
tech sky130A
magscale 1 2
timestamp 1698771642
<< nwell >>
rect 864 676 1684 680
rect 864 672 3592 676
rect -204 650 3592 672
rect -204 608 3304 650
rect -204 578 1896 608
rect -204 204 1044 578
rect 1648 214 1896 578
rect 1904 216 2642 608
rect 1904 214 1974 216
rect 1648 204 1974 214
rect 2306 204 2642 216
rect 842 202 1044 204
rect -34 -598 178 -594
rect 736 -598 1058 -594
rect 1612 -598 1810 -558
rect 2294 -598 3564 -582
rect -34 -604 1183 -598
rect 1612 -604 3564 -598
rect -34 -632 3564 -604
rect -34 -640 6004 -632
rect -34 -1084 6010 -640
rect -34 -1116 6000 -1084
rect 1498 -1126 6000 -1116
rect 2294 -1128 6000 -1126
rect 2294 -1130 3564 -1128
<< nmos >>
rect 556 -2 586 82
rect 756 -2 786 82
rect 256 -478 286 -394
rect 344 -478 374 -394
rect 556 -476 586 -392
rect 756 -476 786 -392
rect 962 -480 992 -396
rect 1162 -482 1192 -398
rect 1364 -480 1394 -396
rect 1564 -482 1594 -398
rect 1990 -482 2020 -398
rect 2086 -482 2116 -398
rect 2182 -482 2212 -398
rect 2404 -482 2434 -398
rect 2500 -482 2530 -398
rect 2596 -482 2626 -398
rect 2692 -482 2722 -398
rect 2788 -482 2818 -398
rect 2884 -482 2914 -398
rect 2980 -482 3010 -398
rect 3076 -482 3106 -398
rect 3172 -482 3202 -398
rect 3380 -482 3410 -398
rect 3476 -482 3506 -398
rect 3572 -482 3602 -398
rect 3668 -482 3698 -398
rect 3764 -482 3794 -398
rect 3860 -482 3890 -398
rect 3956 -482 3986 -398
rect 4052 -482 4082 -398
rect 4148 -482 4178 -398
rect 4244 -482 4274 -398
rect 4340 -482 4370 -398
rect 4436 -482 4466 -398
rect 4532 -482 4562 -398
rect 4628 -482 4658 -398
rect 4724 -482 4754 -398
rect 4820 -482 4850 -398
rect 4916 -482 4946 -398
rect 5012 -482 5042 -398
rect 5108 -482 5138 -398
rect 5204 -482 5234 -398
rect 5300 -482 5330 -398
rect 5396 -482 5426 -398
rect 5492 -482 5522 -398
rect 5588 -482 5618 -398
rect 5684 -482 5714 -398
rect 5780 -482 5810 -398
rect 5876 -482 5906 -398
<< pmos >>
rect 556 266 586 518
rect 756 266 786 518
rect 256 -960 286 -708
rect 344 -960 374 -708
rect 556 -912 586 -660
rect 756 -912 786 -660
rect 962 -918 992 -666
rect 1162 -918 1192 -666
rect 1364 -918 1394 -666
rect 1564 -918 1594 -666
rect 1994 -962 2024 -710
rect 2090 -962 2120 -710
rect 2186 -962 2216 -710
rect 2402 -962 2432 -710
rect 2498 -962 2528 -710
rect 2594 -962 2624 -710
rect 2690 -962 2720 -710
rect 2786 -962 2816 -710
rect 2882 -962 2912 -710
rect 2978 -962 3008 -710
rect 3074 -962 3104 -710
rect 3170 -962 3200 -710
rect 3380 -984 3410 -732
rect 3476 -984 3506 -732
rect 3572 -984 3602 -732
rect 3668 -984 3698 -732
rect 3764 -984 3794 -732
rect 3860 -984 3890 -732
rect 3956 -984 3986 -732
rect 4052 -984 4082 -732
rect 4148 -984 4178 -732
rect 4244 -984 4274 -732
rect 4340 -984 4370 -732
rect 4436 -984 4466 -732
rect 4532 -984 4562 -732
rect 4628 -984 4658 -732
rect 4724 -984 4754 -732
rect 4820 -984 4850 -732
rect 4916 -984 4946 -732
rect 5012 -984 5042 -732
rect 5108 -984 5138 -732
rect 5204 -984 5234 -732
rect 5300 -984 5330 -732
rect 5396 -984 5426 -732
rect 5492 -984 5522 -732
rect 5588 -984 5618 -732
rect 5684 -984 5714 -732
rect 5780 -984 5810 -732
rect 5876 -984 5906 -732
<< ndiff >>
rect 498 70 556 82
rect 498 10 510 70
rect 544 10 556 70
rect 498 -2 556 10
rect 586 70 644 82
rect 586 10 598 70
rect 632 10 644 70
rect 586 -2 644 10
rect 698 70 756 82
rect 698 10 710 70
rect 744 10 756 70
rect 698 -2 756 10
rect 786 70 844 82
rect 786 10 798 70
rect 832 10 844 70
rect 786 -2 844 10
rect 198 -406 256 -394
rect 198 -466 210 -406
rect 244 -466 256 -406
rect 198 -478 256 -466
rect 286 -406 344 -394
rect 286 -466 298 -406
rect 332 -466 344 -406
rect 286 -478 344 -466
rect 374 -406 432 -394
rect 374 -466 386 -406
rect 420 -466 432 -406
rect 374 -478 432 -466
rect 498 -404 556 -392
rect 498 -464 510 -404
rect 544 -464 556 -404
rect 498 -476 556 -464
rect 586 -404 644 -392
rect 586 -464 598 -404
rect 632 -464 644 -404
rect 586 -476 644 -464
rect 698 -404 756 -392
rect 698 -464 710 -404
rect 744 -464 756 -404
rect 698 -476 756 -464
rect 786 -404 844 -392
rect 786 -464 798 -404
rect 832 -464 844 -404
rect 786 -476 844 -464
rect 904 -408 962 -396
rect 904 -468 916 -408
rect 950 -468 962 -408
rect 904 -480 962 -468
rect 992 -408 1050 -396
rect 992 -468 1004 -408
rect 1038 -468 1050 -408
rect 992 -480 1050 -468
rect 1104 -410 1162 -398
rect 1104 -470 1116 -410
rect 1150 -470 1162 -410
rect 1104 -482 1162 -470
rect 1192 -410 1250 -398
rect 1192 -470 1204 -410
rect 1238 -470 1250 -410
rect 1192 -482 1250 -470
rect 1306 -408 1364 -396
rect 1306 -468 1318 -408
rect 1352 -468 1364 -408
rect 1306 -480 1364 -468
rect 1394 -408 1452 -396
rect 1394 -468 1406 -408
rect 1440 -468 1452 -408
rect 1394 -480 1452 -468
rect 1506 -410 1564 -398
rect 1506 -470 1518 -410
rect 1552 -470 1564 -410
rect 1506 -482 1564 -470
rect 1594 -410 1652 -398
rect 1594 -470 1606 -410
rect 1640 -470 1652 -410
rect 1594 -482 1652 -470
rect 1928 -410 1990 -398
rect 1928 -470 1940 -410
rect 1974 -470 1990 -410
rect 1928 -482 1990 -470
rect 2020 -410 2086 -398
rect 2020 -470 2036 -410
rect 2070 -470 2086 -410
rect 2020 -482 2086 -470
rect 2116 -410 2182 -398
rect 2116 -470 2132 -410
rect 2166 -470 2182 -410
rect 2116 -482 2182 -470
rect 2212 -410 2274 -398
rect 2212 -470 2228 -410
rect 2262 -470 2274 -410
rect 2212 -482 2274 -470
rect 2342 -410 2404 -398
rect 2342 -470 2354 -410
rect 2388 -470 2404 -410
rect 2342 -482 2404 -470
rect 2434 -410 2500 -398
rect 2434 -470 2450 -410
rect 2484 -470 2500 -410
rect 2434 -482 2500 -470
rect 2530 -410 2596 -398
rect 2530 -470 2546 -410
rect 2580 -470 2596 -410
rect 2530 -482 2596 -470
rect 2626 -410 2692 -398
rect 2626 -470 2642 -410
rect 2676 -470 2692 -410
rect 2626 -482 2692 -470
rect 2722 -410 2788 -398
rect 2722 -470 2738 -410
rect 2772 -470 2788 -410
rect 2722 -482 2788 -470
rect 2818 -410 2884 -398
rect 2818 -470 2834 -410
rect 2868 -470 2884 -410
rect 2818 -482 2884 -470
rect 2914 -410 2980 -398
rect 2914 -470 2930 -410
rect 2964 -470 2980 -410
rect 2914 -482 2980 -470
rect 3010 -410 3076 -398
rect 3010 -470 3026 -410
rect 3060 -470 3076 -410
rect 3010 -482 3076 -470
rect 3106 -410 3172 -398
rect 3106 -470 3122 -410
rect 3156 -470 3172 -410
rect 3106 -482 3172 -470
rect 3202 -410 3264 -398
rect 3202 -470 3218 -410
rect 3252 -470 3264 -410
rect 3202 -482 3264 -470
rect 3318 -410 3380 -398
rect 3318 -470 3330 -410
rect 3364 -470 3380 -410
rect 3318 -482 3380 -470
rect 3410 -410 3476 -398
rect 3410 -470 3426 -410
rect 3460 -470 3476 -410
rect 3410 -482 3476 -470
rect 3506 -410 3572 -398
rect 3506 -470 3522 -410
rect 3556 -470 3572 -410
rect 3506 -482 3572 -470
rect 3602 -410 3668 -398
rect 3602 -470 3618 -410
rect 3652 -470 3668 -410
rect 3602 -482 3668 -470
rect 3698 -410 3764 -398
rect 3698 -470 3714 -410
rect 3748 -470 3764 -410
rect 3698 -482 3764 -470
rect 3794 -410 3860 -398
rect 3794 -470 3810 -410
rect 3844 -470 3860 -410
rect 3794 -482 3860 -470
rect 3890 -410 3956 -398
rect 3890 -470 3906 -410
rect 3940 -470 3956 -410
rect 3890 -482 3956 -470
rect 3986 -410 4052 -398
rect 3986 -470 4002 -410
rect 4036 -470 4052 -410
rect 3986 -482 4052 -470
rect 4082 -410 4148 -398
rect 4082 -470 4098 -410
rect 4132 -470 4148 -410
rect 4082 -482 4148 -470
rect 4178 -410 4244 -398
rect 4178 -470 4194 -410
rect 4228 -470 4244 -410
rect 4178 -482 4244 -470
rect 4274 -410 4340 -398
rect 4274 -470 4290 -410
rect 4324 -470 4340 -410
rect 4274 -482 4340 -470
rect 4370 -410 4436 -398
rect 4370 -470 4386 -410
rect 4420 -470 4436 -410
rect 4370 -482 4436 -470
rect 4466 -410 4532 -398
rect 4466 -470 4482 -410
rect 4516 -470 4532 -410
rect 4466 -482 4532 -470
rect 4562 -410 4628 -398
rect 4562 -470 4578 -410
rect 4612 -470 4628 -410
rect 4562 -482 4628 -470
rect 4658 -410 4724 -398
rect 4658 -470 4674 -410
rect 4708 -470 4724 -410
rect 4658 -482 4724 -470
rect 4754 -410 4820 -398
rect 4754 -470 4770 -410
rect 4804 -470 4820 -410
rect 4754 -482 4820 -470
rect 4850 -410 4916 -398
rect 4850 -470 4866 -410
rect 4900 -470 4916 -410
rect 4850 -482 4916 -470
rect 4946 -410 5012 -398
rect 4946 -470 4962 -410
rect 4996 -470 5012 -410
rect 4946 -482 5012 -470
rect 5042 -410 5108 -398
rect 5042 -470 5058 -410
rect 5092 -470 5108 -410
rect 5042 -482 5108 -470
rect 5138 -410 5204 -398
rect 5138 -470 5154 -410
rect 5188 -470 5204 -410
rect 5138 -482 5204 -470
rect 5234 -410 5300 -398
rect 5234 -470 5250 -410
rect 5284 -470 5300 -410
rect 5234 -482 5300 -470
rect 5330 -410 5396 -398
rect 5330 -470 5346 -410
rect 5380 -470 5396 -410
rect 5330 -482 5396 -470
rect 5426 -410 5492 -398
rect 5426 -470 5442 -410
rect 5476 -470 5492 -410
rect 5426 -482 5492 -470
rect 5522 -410 5588 -398
rect 5522 -470 5538 -410
rect 5572 -470 5588 -410
rect 5522 -482 5588 -470
rect 5618 -410 5684 -398
rect 5618 -470 5634 -410
rect 5668 -470 5684 -410
rect 5618 -482 5684 -470
rect 5714 -410 5780 -398
rect 5714 -470 5730 -410
rect 5764 -470 5780 -410
rect 5714 -482 5780 -470
rect 5810 -410 5876 -398
rect 5810 -470 5826 -410
rect 5860 -470 5876 -410
rect 5810 -482 5876 -470
rect 5906 -410 5968 -398
rect 5906 -470 5922 -410
rect 5956 -470 5968 -410
rect 5906 -482 5968 -470
<< pdiff >>
rect 498 506 556 518
rect 498 278 510 506
rect 544 278 556 506
rect 498 266 556 278
rect 586 506 644 518
rect 586 278 598 506
rect 632 278 644 506
rect 586 266 644 278
rect 698 506 756 518
rect 698 278 710 506
rect 744 278 756 506
rect 698 266 756 278
rect 786 506 844 518
rect 786 278 798 506
rect 832 278 844 506
rect 786 266 844 278
rect 498 -672 556 -660
rect 198 -720 256 -708
rect 198 -948 210 -720
rect 244 -948 256 -720
rect 198 -960 256 -948
rect 286 -720 344 -708
rect 286 -948 298 -720
rect 332 -948 344 -720
rect 286 -960 344 -948
rect 374 -720 432 -708
rect 374 -948 386 -720
rect 420 -948 432 -720
rect 498 -900 510 -672
rect 544 -900 556 -672
rect 498 -912 556 -900
rect 586 -672 644 -660
rect 586 -900 598 -672
rect 632 -900 644 -672
rect 586 -912 644 -900
rect 698 -672 756 -660
rect 698 -900 710 -672
rect 744 -900 756 -672
rect 698 -912 756 -900
rect 786 -672 844 -660
rect 786 -900 798 -672
rect 832 -900 844 -672
rect 786 -912 844 -900
rect 904 -678 962 -666
rect 904 -906 916 -678
rect 950 -906 962 -678
rect 374 -960 432 -948
rect 904 -918 962 -906
rect 992 -678 1050 -666
rect 992 -906 1004 -678
rect 1038 -906 1050 -678
rect 992 -918 1050 -906
rect 1104 -678 1162 -666
rect 1104 -906 1116 -678
rect 1150 -906 1162 -678
rect 1104 -918 1162 -906
rect 1192 -678 1250 -666
rect 1192 -906 1204 -678
rect 1238 -906 1250 -678
rect 1192 -918 1250 -906
rect 1306 -678 1364 -666
rect 1306 -906 1318 -678
rect 1352 -906 1364 -678
rect 1306 -918 1364 -906
rect 1394 -678 1452 -666
rect 1394 -906 1406 -678
rect 1440 -906 1452 -678
rect 1394 -918 1452 -906
rect 1506 -678 1564 -666
rect 1506 -906 1518 -678
rect 1552 -906 1564 -678
rect 1506 -918 1564 -906
rect 1594 -678 1652 -666
rect 1594 -906 1606 -678
rect 1640 -906 1652 -678
rect 1594 -918 1652 -906
rect 1932 -722 1994 -710
rect 1932 -950 1944 -722
rect 1978 -950 1994 -722
rect 1932 -962 1994 -950
rect 2024 -722 2090 -710
rect 2024 -950 2040 -722
rect 2074 -950 2090 -722
rect 2024 -962 2090 -950
rect 2120 -722 2186 -710
rect 2120 -950 2136 -722
rect 2170 -950 2186 -722
rect 2120 -962 2186 -950
rect 2216 -722 2278 -710
rect 2216 -950 2232 -722
rect 2266 -950 2278 -722
rect 2216 -962 2278 -950
rect 2340 -722 2402 -710
rect 2340 -950 2352 -722
rect 2386 -950 2402 -722
rect 2340 -962 2402 -950
rect 2432 -722 2498 -710
rect 2432 -950 2448 -722
rect 2482 -950 2498 -722
rect 2432 -962 2498 -950
rect 2528 -722 2594 -710
rect 2528 -950 2544 -722
rect 2578 -950 2594 -722
rect 2528 -962 2594 -950
rect 2624 -722 2690 -710
rect 2624 -950 2640 -722
rect 2674 -950 2690 -722
rect 2624 -962 2690 -950
rect 2720 -722 2786 -710
rect 2720 -950 2736 -722
rect 2770 -950 2786 -722
rect 2720 -962 2786 -950
rect 2816 -722 2882 -710
rect 2816 -950 2832 -722
rect 2866 -950 2882 -722
rect 2816 -962 2882 -950
rect 2912 -722 2978 -710
rect 2912 -950 2928 -722
rect 2962 -950 2978 -722
rect 2912 -962 2978 -950
rect 3008 -722 3074 -710
rect 3008 -950 3024 -722
rect 3058 -950 3074 -722
rect 3008 -962 3074 -950
rect 3104 -722 3170 -710
rect 3104 -950 3120 -722
rect 3154 -950 3170 -722
rect 3104 -962 3170 -950
rect 3200 -722 3262 -710
rect 3200 -950 3216 -722
rect 3250 -950 3262 -722
rect 3200 -962 3262 -950
rect 3318 -744 3380 -732
rect 3318 -972 3330 -744
rect 3364 -972 3380 -744
rect 3318 -984 3380 -972
rect 3410 -744 3476 -732
rect 3410 -972 3426 -744
rect 3460 -972 3476 -744
rect 3410 -984 3476 -972
rect 3506 -744 3572 -732
rect 3506 -972 3522 -744
rect 3556 -972 3572 -744
rect 3506 -984 3572 -972
rect 3602 -744 3668 -732
rect 3602 -972 3618 -744
rect 3652 -972 3668 -744
rect 3602 -984 3668 -972
rect 3698 -744 3764 -732
rect 3698 -972 3714 -744
rect 3748 -972 3764 -744
rect 3698 -984 3764 -972
rect 3794 -744 3860 -732
rect 3794 -972 3810 -744
rect 3844 -972 3860 -744
rect 3794 -984 3860 -972
rect 3890 -744 3956 -732
rect 3890 -972 3906 -744
rect 3940 -972 3956 -744
rect 3890 -984 3956 -972
rect 3986 -744 4052 -732
rect 3986 -972 4002 -744
rect 4036 -972 4052 -744
rect 3986 -984 4052 -972
rect 4082 -744 4148 -732
rect 4082 -972 4098 -744
rect 4132 -972 4148 -744
rect 4082 -984 4148 -972
rect 4178 -744 4244 -732
rect 4178 -972 4194 -744
rect 4228 -972 4244 -744
rect 4178 -984 4244 -972
rect 4274 -744 4340 -732
rect 4274 -972 4290 -744
rect 4324 -972 4340 -744
rect 4274 -984 4340 -972
rect 4370 -744 4436 -732
rect 4370 -972 4386 -744
rect 4420 -972 4436 -744
rect 4370 -984 4436 -972
rect 4466 -744 4532 -732
rect 4466 -972 4482 -744
rect 4516 -972 4532 -744
rect 4466 -984 4532 -972
rect 4562 -744 4628 -732
rect 4562 -972 4578 -744
rect 4612 -972 4628 -744
rect 4562 -984 4628 -972
rect 4658 -744 4724 -732
rect 4658 -972 4674 -744
rect 4708 -972 4724 -744
rect 4658 -984 4724 -972
rect 4754 -744 4820 -732
rect 4754 -972 4770 -744
rect 4804 -972 4820 -744
rect 4754 -984 4820 -972
rect 4850 -744 4916 -732
rect 4850 -972 4866 -744
rect 4900 -972 4916 -744
rect 4850 -984 4916 -972
rect 4946 -744 5012 -732
rect 4946 -972 4962 -744
rect 4996 -972 5012 -744
rect 4946 -984 5012 -972
rect 5042 -744 5108 -732
rect 5042 -972 5058 -744
rect 5092 -972 5108 -744
rect 5042 -984 5108 -972
rect 5138 -744 5204 -732
rect 5138 -972 5154 -744
rect 5188 -972 5204 -744
rect 5138 -984 5204 -972
rect 5234 -744 5300 -732
rect 5234 -972 5250 -744
rect 5284 -972 5300 -744
rect 5234 -984 5300 -972
rect 5330 -744 5396 -732
rect 5330 -972 5346 -744
rect 5380 -972 5396 -744
rect 5330 -984 5396 -972
rect 5426 -744 5492 -732
rect 5426 -972 5442 -744
rect 5476 -972 5492 -744
rect 5426 -984 5492 -972
rect 5522 -744 5588 -732
rect 5522 -972 5538 -744
rect 5572 -972 5588 -744
rect 5522 -984 5588 -972
rect 5618 -744 5684 -732
rect 5618 -972 5634 -744
rect 5668 -972 5684 -744
rect 5618 -984 5684 -972
rect 5714 -744 5780 -732
rect 5714 -972 5730 -744
rect 5764 -972 5780 -744
rect 5714 -984 5780 -972
rect 5810 -744 5876 -732
rect 5810 -972 5826 -744
rect 5860 -972 5876 -744
rect 5810 -984 5876 -972
rect 5906 -744 5968 -732
rect 5906 -972 5922 -744
rect 5956 -972 5968 -744
rect 5906 -984 5968 -972
<< ndiffc >>
rect 510 10 544 70
rect 598 10 632 70
rect 710 10 744 70
rect 798 10 832 70
rect 210 -466 244 -406
rect 298 -466 332 -406
rect 386 -466 420 -406
rect 510 -464 544 -404
rect 598 -464 632 -404
rect 710 -464 744 -404
rect 798 -464 832 -404
rect 916 -468 950 -408
rect 1004 -468 1038 -408
rect 1116 -470 1150 -410
rect 1204 -470 1238 -410
rect 1318 -468 1352 -408
rect 1406 -468 1440 -408
rect 1518 -470 1552 -410
rect 1606 -470 1640 -410
rect 1940 -470 1974 -410
rect 2036 -470 2070 -410
rect 2132 -470 2166 -410
rect 2228 -470 2262 -410
rect 2354 -470 2388 -410
rect 2450 -470 2484 -410
rect 2546 -470 2580 -410
rect 2642 -470 2676 -410
rect 2738 -470 2772 -410
rect 2834 -470 2868 -410
rect 2930 -470 2964 -410
rect 3026 -470 3060 -410
rect 3122 -470 3156 -410
rect 3218 -470 3252 -410
rect 3330 -470 3364 -410
rect 3426 -470 3460 -410
rect 3522 -470 3556 -410
rect 3618 -470 3652 -410
rect 3714 -470 3748 -410
rect 3810 -470 3844 -410
rect 3906 -470 3940 -410
rect 4002 -470 4036 -410
rect 4098 -470 4132 -410
rect 4194 -470 4228 -410
rect 4290 -470 4324 -410
rect 4386 -470 4420 -410
rect 4482 -470 4516 -410
rect 4578 -470 4612 -410
rect 4674 -470 4708 -410
rect 4770 -470 4804 -410
rect 4866 -470 4900 -410
rect 4962 -470 4996 -410
rect 5058 -470 5092 -410
rect 5154 -470 5188 -410
rect 5250 -470 5284 -410
rect 5346 -470 5380 -410
rect 5442 -470 5476 -410
rect 5538 -470 5572 -410
rect 5634 -470 5668 -410
rect 5730 -470 5764 -410
rect 5826 -470 5860 -410
rect 5922 -470 5956 -410
<< pdiffc >>
rect 510 278 544 506
rect 598 278 632 506
rect 710 278 744 506
rect 798 278 832 506
rect 210 -948 244 -720
rect 298 -948 332 -720
rect 386 -948 420 -720
rect 510 -900 544 -672
rect 598 -900 632 -672
rect 710 -900 744 -672
rect 798 -900 832 -672
rect 916 -906 950 -678
rect 1004 -906 1038 -678
rect 1116 -906 1150 -678
rect 1204 -906 1238 -678
rect 1318 -906 1352 -678
rect 1406 -906 1440 -678
rect 1518 -906 1552 -678
rect 1606 -906 1640 -678
rect 1944 -950 1978 -722
rect 2040 -950 2074 -722
rect 2136 -950 2170 -722
rect 2232 -950 2266 -722
rect 2352 -950 2386 -722
rect 2448 -950 2482 -722
rect 2544 -950 2578 -722
rect 2640 -950 2674 -722
rect 2736 -950 2770 -722
rect 2832 -950 2866 -722
rect 2928 -950 2962 -722
rect 3024 -950 3058 -722
rect 3120 -950 3154 -722
rect 3216 -950 3250 -722
rect 3330 -972 3364 -744
rect 3426 -972 3460 -744
rect 3522 -972 3556 -744
rect 3618 -972 3652 -744
rect 3714 -972 3748 -744
rect 3810 -972 3844 -744
rect 3906 -972 3940 -744
rect 4002 -972 4036 -744
rect 4098 -972 4132 -744
rect 4194 -972 4228 -744
rect 4290 -972 4324 -744
rect 4386 -972 4420 -744
rect 4482 -972 4516 -744
rect 4578 -972 4612 -744
rect 4674 -972 4708 -744
rect 4770 -972 4804 -744
rect 4866 -972 4900 -744
rect 4962 -972 4996 -744
rect 5058 -972 5092 -744
rect 5154 -972 5188 -744
rect 5250 -972 5284 -744
rect 5346 -972 5380 -744
rect 5442 -972 5476 -744
rect 5538 -972 5572 -744
rect 5634 -972 5668 -744
rect 5730 -972 5764 -744
rect 5826 -972 5860 -744
rect 5922 -972 5956 -744
<< psubdiff >>
rect 24 -412 112 -394
rect 24 -460 48 -412
rect 86 -460 112 -412
rect 24 -480 112 -460
<< nsubdiff >>
rect -162 578 -76 606
rect -162 290 -138 578
rect -100 290 -76 578
rect -162 258 -76 290
rect 2 -732 76 -706
rect 2 -928 22 -732
rect 56 -928 76 -732
rect 2 -954 76 -928
<< psubdiffcont >>
rect 48 -460 86 -412
<< nsubdiffcont >>
rect -138 290 -100 578
rect 22 -928 56 -732
<< poly >>
rect 618 646 792 654
rect 618 638 794 646
rect 618 604 638 638
rect 778 604 794 638
rect 618 592 794 604
rect 1994 612 2216 648
rect 618 588 792 592
rect 556 518 586 544
rect 756 518 786 588
rect 1994 570 2024 612
rect 2186 576 2216 612
rect 2402 614 3200 648
rect 2402 572 2432 614
rect 2594 572 2624 614
rect 2786 570 2816 614
rect 2978 570 3008 614
rect 3170 570 3200 614
rect 56 198 86 266
rect 256 200 286 290
rect -40 196 88 198
rect -44 180 88 196
rect -44 136 -28 180
rect 72 136 88 180
rect -44 122 88 136
rect 134 180 286 200
rect 134 140 146 180
rect 272 140 286 180
rect 134 122 286 140
rect -44 120 86 122
rect 136 120 286 122
rect 56 100 86 120
rect 256 104 286 120
rect 344 102 374 294
rect 556 198 586 266
rect 416 180 586 198
rect 416 140 440 180
rect 570 140 586 180
rect 416 120 586 140
rect 556 82 586 120
rect 756 82 786 266
rect 956 220 986 260
rect 1156 226 1186 266
rect 1358 230 1388 268
rect 1992 266 2026 278
rect 2090 266 2120 314
rect 2498 268 2528 312
rect 2690 268 2720 310
rect 2882 268 2912 312
rect 3074 268 3104 312
rect 1558 230 1588 262
rect 1976 234 2234 266
rect 2384 234 3201 268
rect 1992 233 2026 234
rect 1990 232 2026 233
rect 832 206 986 220
rect 832 144 848 206
rect 946 144 986 206
rect 832 132 986 144
rect 956 96 986 132
rect 1028 212 1188 226
rect 1028 138 1046 212
rect 1144 138 1188 212
rect 1028 120 1188 138
rect 1230 214 1388 230
rect 1230 140 1246 214
rect 1344 140 1388 214
rect 1230 122 1388 140
rect 1430 214 1588 230
rect 1430 140 1446 214
rect 1544 140 1588 214
rect 1976 216 2026 232
rect 1976 192 2024 216
rect 2384 204 2436 234
rect 1430 122 1588 140
rect 1648 176 2024 192
rect 1648 138 1664 176
rect 1926 158 2024 176
rect 2280 190 2436 204
rect 1926 138 2212 158
rect 2280 148 2298 190
rect 2370 158 2436 190
rect 3246 166 3400 182
rect 2370 148 3202 158
rect 2280 138 3202 148
rect 1648 126 2212 138
rect 1948 124 2212 126
rect 1156 102 1186 120
rect 1358 104 1388 122
rect 1558 98 1588 122
rect 1990 110 2022 124
rect 1990 94 2020 110
rect 2182 94 2212 124
rect 2404 126 3202 138
rect 2404 86 2434 126
rect 2596 86 2626 126
rect 2788 88 2818 126
rect 2980 88 3010 126
rect 3172 94 3202 126
rect 3246 130 3264 166
rect 3384 130 3400 166
rect 3246 124 3400 130
rect 3246 118 3398 124
rect 3175 93 3201 94
rect 338 -74 374 -20
rect 556 -28 586 -2
rect 756 -28 786 -2
rect 2086 -36 2116 0
rect 2500 -36 2530 -2
rect 2692 -36 2722 0
rect 2884 -36 2914 4
rect 3076 -36 3106 4
rect 1972 -70 2230 -36
rect 2387 -70 3220 -36
rect 2500 -72 2530 -70
rect 338 -86 792 -74
rect 338 -122 354 -86
rect 770 -122 792 -86
rect 338 -132 792 -122
rect 344 -248 798 -236
rect 344 -302 360 -248
rect 780 -302 798 -248
rect 344 -312 798 -302
rect 256 -394 286 -368
rect 344 -394 374 -312
rect 1972 -326 2038 -310
rect 2164 -326 2230 -310
rect 1972 -360 1988 -326
rect 2022 -360 2180 -326
rect 2214 -360 2230 -326
rect 556 -392 586 -366
rect 756 -392 786 -366
rect 962 -396 992 -370
rect 256 -516 286 -478
rect -56 -534 286 -516
rect -56 -576 -40 -534
rect 272 -576 286 -534
rect -56 -592 286 -576
rect 210 -594 286 -592
rect 256 -708 286 -594
rect 344 -708 374 -478
rect 556 -514 586 -476
rect 420 -534 586 -514
rect 420 -576 432 -534
rect 570 -576 586 -534
rect 420 -594 586 -576
rect 556 -660 586 -594
rect 756 -660 786 -476
rect 1162 -398 1192 -372
rect 1364 -396 1394 -370
rect 962 -518 992 -480
rect 1564 -398 1594 -372
rect 1972 -376 2038 -360
rect 1990 -398 2020 -376
rect 2086 -398 2116 -360
rect 2164 -376 2230 -360
rect 2386 -326 2452 -310
rect 2500 -326 2530 -324
rect 2578 -326 2644 -310
rect 2770 -326 2836 -310
rect 2962 -326 3028 -310
rect 3154 -326 3220 -310
rect 3362 -326 3428 -310
rect 3554 -326 3620 -310
rect 3746 -326 3812 -310
rect 3938 -326 4004 -310
rect 4130 -326 4196 -310
rect 4322 -326 4388 -310
rect 4514 -326 4580 -310
rect 4706 -326 4772 -310
rect 4898 -326 4964 -310
rect 5090 -326 5156 -310
rect 5282 -326 5348 -310
rect 5474 -326 5540 -310
rect 5666 -326 5732 -310
rect 5858 -326 5924 -310
rect 2386 -360 2402 -326
rect 2436 -360 2594 -326
rect 2628 -360 2786 -326
rect 2820 -360 2978 -326
rect 3012 -360 3170 -326
rect 3204 -360 3220 -326
rect 3361 -360 3378 -326
rect 3412 -360 3570 -326
rect 3604 -360 3762 -326
rect 3796 -360 3954 -326
rect 3988 -360 4146 -326
rect 4180 -360 4338 -326
rect 4372 -360 4530 -326
rect 4564 -360 4722 -326
rect 4756 -360 4914 -326
rect 4948 -360 5106 -326
rect 5140 -360 5298 -326
rect 5332 -360 5490 -326
rect 5524 -360 5682 -326
rect 5716 -360 5874 -326
rect 5908 -360 5924 -326
rect 2386 -376 2452 -360
rect 2182 -398 2212 -376
rect 2404 -398 2434 -376
rect 2500 -398 2530 -360
rect 2578 -376 2644 -360
rect 2596 -398 2626 -376
rect 2692 -398 2722 -360
rect 2770 -376 2836 -360
rect 2788 -398 2818 -376
rect 2884 -398 2914 -360
rect 2962 -376 3028 -360
rect 2980 -398 3010 -376
rect 3076 -398 3106 -360
rect 3154 -376 3220 -360
rect 3362 -376 3428 -360
rect 3172 -398 3202 -376
rect 3380 -398 3410 -376
rect 3476 -398 3506 -360
rect 3554 -376 3620 -360
rect 3572 -398 3602 -376
rect 3668 -398 3698 -360
rect 3746 -376 3812 -360
rect 3764 -398 3794 -376
rect 3860 -398 3890 -360
rect 3938 -376 4004 -360
rect 3956 -398 3986 -376
rect 4052 -398 4082 -360
rect 4130 -376 4196 -360
rect 4148 -398 4178 -376
rect 4244 -398 4274 -360
rect 4322 -376 4388 -360
rect 4340 -398 4370 -376
rect 4436 -398 4466 -360
rect 4514 -376 4580 -360
rect 4532 -398 4562 -376
rect 4628 -398 4658 -360
rect 4706 -376 4772 -360
rect 4724 -398 4754 -376
rect 4820 -398 4850 -360
rect 4898 -376 4964 -360
rect 4916 -398 4946 -376
rect 5012 -398 5042 -360
rect 5090 -376 5156 -360
rect 5108 -398 5138 -376
rect 5204 -398 5234 -360
rect 5282 -376 5348 -360
rect 5300 -398 5330 -376
rect 5396 -398 5426 -360
rect 5474 -376 5540 -360
rect 5492 -398 5522 -376
rect 5588 -398 5618 -360
rect 5666 -376 5732 -360
rect 5684 -398 5714 -376
rect 5780 -398 5810 -360
rect 5858 -376 5924 -360
rect 5876 -398 5906 -376
rect 1162 -518 1192 -482
rect 828 -530 992 -518
rect 828 -568 844 -530
rect 948 -568 992 -530
rect 828 -580 992 -568
rect 962 -666 992 -580
rect 1034 -536 1194 -518
rect 1364 -520 1394 -480
rect 1564 -520 1594 -482
rect 1990 -506 2020 -482
rect 2086 -504 2116 -482
rect 1034 -610 1052 -536
rect 1150 -610 1194 -536
rect 1034 -624 1194 -610
rect 1236 -538 1394 -520
rect 1236 -612 1252 -538
rect 1350 -612 1394 -538
rect 1162 -666 1192 -624
rect 1236 -628 1394 -612
rect 1436 -538 1594 -520
rect 1436 -612 1452 -538
rect 1550 -612 1594 -538
rect 1678 -518 2020 -506
rect 1678 -576 1698 -518
rect 1858 -520 2020 -518
rect 2068 -520 2134 -504
rect 2182 -520 2212 -482
rect 1858 -554 2084 -520
rect 2118 -554 2212 -520
rect 2404 -522 2434 -482
rect 2500 -504 2530 -482
rect 2482 -520 2548 -504
rect 2482 -522 2498 -520
rect 2404 -536 2498 -522
rect 2278 -548 2498 -536
rect 1858 -576 2024 -554
rect 2068 -570 2134 -554
rect 1678 -588 2024 -576
rect 1436 -628 1594 -612
rect 1364 -666 1394 -628
rect 1564 -666 1594 -628
rect 1976 -612 2024 -588
rect 2278 -582 2296 -548
rect 2392 -554 2498 -548
rect 2532 -522 2548 -520
rect 2596 -522 2626 -482
rect 2692 -504 2722 -482
rect 2674 -520 2740 -504
rect 2674 -522 2690 -520
rect 2532 -554 2690 -522
rect 2724 -522 2740 -520
rect 2788 -522 2818 -482
rect 2884 -504 2914 -482
rect 2866 -520 2932 -504
rect 2866 -522 2882 -520
rect 2724 -554 2882 -522
rect 2916 -522 2932 -520
rect 2980 -522 3010 -482
rect 3076 -504 3106 -482
rect 3058 -520 3124 -504
rect 3058 -522 3074 -520
rect 2916 -554 3074 -522
rect 3108 -522 3124 -520
rect 3172 -522 3202 -482
rect 3380 -520 3410 -482
rect 3476 -504 3506 -482
rect 3108 -554 3202 -522
rect 3252 -521 3410 -520
rect 3458 -520 3524 -504
rect 3458 -521 3474 -520
rect 3252 -532 3474 -521
rect 2392 -582 2436 -554
rect 2482 -570 2548 -554
rect 2674 -570 2740 -554
rect 2866 -570 2932 -554
rect 3058 -570 3124 -554
rect 3252 -570 3270 -532
rect 3374 -554 3474 -532
rect 3508 -521 3524 -520
rect 3572 -521 3602 -482
rect 3668 -504 3698 -482
rect 3650 -520 3716 -504
rect 3650 -521 3666 -520
rect 3508 -554 3666 -521
rect 3700 -521 3716 -520
rect 3764 -521 3794 -482
rect 3860 -504 3890 -482
rect 3842 -520 3908 -504
rect 3842 -521 3858 -520
rect 3700 -554 3858 -521
rect 3892 -521 3908 -520
rect 3956 -521 3986 -482
rect 4052 -504 4082 -482
rect 4034 -520 4100 -504
rect 4034 -521 4050 -520
rect 3892 -554 4050 -521
rect 4084 -521 4100 -520
rect 4148 -521 4178 -482
rect 4244 -504 4274 -482
rect 4226 -520 4292 -504
rect 4226 -521 4242 -520
rect 4084 -554 4242 -521
rect 4276 -521 4292 -520
rect 4340 -521 4370 -482
rect 4436 -504 4466 -482
rect 4418 -520 4484 -504
rect 4418 -521 4434 -520
rect 4276 -554 4434 -521
rect 4468 -521 4484 -520
rect 4532 -521 4562 -482
rect 4628 -504 4658 -482
rect 4610 -520 4676 -504
rect 4610 -521 4626 -520
rect 4468 -554 4626 -521
rect 4660 -521 4676 -520
rect 4724 -521 4754 -482
rect 4820 -504 4850 -482
rect 4802 -520 4868 -504
rect 4802 -521 4818 -520
rect 4660 -554 4818 -521
rect 4852 -521 4868 -520
rect 4916 -521 4946 -482
rect 5012 -504 5042 -482
rect 4994 -520 5060 -504
rect 4994 -521 5010 -520
rect 4852 -554 5010 -521
rect 5044 -521 5060 -520
rect 5108 -521 5138 -482
rect 5204 -504 5234 -482
rect 5186 -520 5252 -504
rect 5186 -521 5202 -520
rect 5044 -554 5202 -521
rect 5236 -521 5252 -520
rect 5300 -521 5330 -482
rect 5396 -504 5426 -482
rect 5378 -520 5444 -504
rect 5378 -521 5394 -520
rect 5236 -554 5394 -521
rect 5428 -521 5444 -520
rect 5492 -521 5522 -482
rect 5588 -504 5618 -482
rect 5570 -520 5636 -504
rect 5570 -521 5586 -520
rect 5428 -554 5586 -521
rect 5620 -521 5636 -520
rect 5684 -521 5714 -482
rect 5780 -504 5810 -482
rect 5762 -520 5828 -504
rect 5762 -521 5778 -520
rect 5620 -554 5778 -521
rect 5812 -521 5828 -520
rect 5876 -521 5906 -482
rect 5812 -554 5909 -521
rect 3374 -555 5909 -554
rect 3374 -570 3410 -555
rect 3458 -570 3524 -555
rect 3650 -570 3716 -555
rect 3842 -570 3908 -555
rect 3956 -556 3986 -555
rect 4034 -570 4100 -555
rect 4226 -570 4292 -555
rect 4418 -570 4484 -555
rect 4610 -570 4676 -555
rect 4802 -570 4868 -555
rect 4994 -570 5060 -555
rect 5186 -570 5252 -555
rect 5378 -570 5444 -555
rect 5492 -556 5522 -555
rect 5570 -570 5636 -555
rect 5684 -556 5714 -555
rect 5762 -570 5828 -555
rect 3252 -582 3410 -570
rect 5875 -578 5909 -555
rect 2278 -594 2436 -582
rect 1976 -613 2026 -612
rect 2384 -613 2436 -594
rect 1976 -629 2042 -613
rect 1976 -663 1992 -629
rect 2026 -630 2042 -629
rect 2168 -629 2234 -613
rect 2168 -630 2184 -629
rect 2026 -662 2184 -630
rect 2026 -663 2042 -662
rect 556 -938 586 -912
rect 256 -986 286 -960
rect 344 -986 374 -960
rect 756 -986 786 -912
rect 1976 -679 2042 -663
rect 1994 -710 2024 -679
rect 2090 -710 2120 -662
rect 2168 -663 2184 -662
rect 2218 -663 2234 -629
rect 2168 -679 2234 -663
rect 2384 -629 2450 -613
rect 2384 -663 2400 -629
rect 2434 -630 2450 -629
rect 2576 -629 2642 -613
rect 2576 -630 2592 -629
rect 2434 -663 2592 -630
rect 2626 -630 2642 -629
rect 2768 -629 2834 -613
rect 2768 -630 2784 -629
rect 2626 -663 2784 -630
rect 2818 -630 2834 -629
rect 2960 -629 3026 -613
rect 2960 -630 2976 -629
rect 2818 -663 2976 -630
rect 3010 -630 3026 -629
rect 3152 -629 3218 -613
rect 3152 -630 3168 -629
rect 3010 -663 3168 -630
rect 3202 -663 3218 -629
rect 3380 -635 3410 -582
rect 5876 -635 5906 -578
rect 3362 -651 3428 -635
rect 3362 -658 3378 -651
rect 2384 -664 3218 -663
rect 2384 -679 2450 -664
rect 2186 -710 2216 -679
rect 2402 -710 2432 -679
rect 2498 -710 2528 -664
rect 2576 -679 2642 -664
rect 2594 -710 2624 -679
rect 2690 -710 2720 -664
rect 2768 -679 2834 -664
rect 2786 -710 2816 -679
rect 2882 -710 2912 -664
rect 2960 -679 3026 -664
rect 2978 -710 3008 -679
rect 3074 -710 3104 -664
rect 3152 -679 3218 -664
rect 3170 -710 3200 -679
rect 3360 -685 3378 -658
rect 3412 -658 3428 -651
rect 3554 -651 3620 -635
rect 3554 -658 3570 -651
rect 3412 -685 3570 -658
rect 3604 -658 3620 -651
rect 3746 -651 3812 -635
rect 3746 -658 3762 -651
rect 3604 -685 3762 -658
rect 3796 -658 3812 -651
rect 3938 -651 4004 -635
rect 3938 -658 3954 -651
rect 3796 -685 3954 -658
rect 3988 -658 4004 -651
rect 4130 -651 4196 -635
rect 4130 -658 4146 -651
rect 3988 -685 4146 -658
rect 4180 -658 4196 -651
rect 4322 -651 4388 -635
rect 4322 -658 4338 -651
rect 4180 -685 4338 -658
rect 4372 -658 4388 -651
rect 4514 -651 4580 -635
rect 4514 -658 4530 -651
rect 4372 -685 4530 -658
rect 4564 -658 4580 -651
rect 4706 -651 4772 -635
rect 4706 -658 4722 -651
rect 4564 -685 4722 -658
rect 4756 -658 4772 -651
rect 4898 -651 4964 -635
rect 4898 -658 4914 -651
rect 4756 -685 4914 -658
rect 4948 -658 4964 -651
rect 5090 -651 5156 -635
rect 5090 -658 5106 -651
rect 4948 -685 5106 -658
rect 5140 -658 5156 -651
rect 5282 -651 5348 -635
rect 5282 -658 5298 -651
rect 5140 -685 5298 -658
rect 5332 -658 5348 -651
rect 5474 -651 5540 -635
rect 5474 -658 5490 -651
rect 5332 -685 5490 -658
rect 5524 -658 5540 -651
rect 5666 -651 5732 -635
rect 5666 -658 5682 -651
rect 5524 -685 5682 -658
rect 5716 -658 5732 -651
rect 5858 -651 5924 -635
rect 5858 -658 5874 -651
rect 5716 -685 5874 -658
rect 5908 -685 5924 -651
rect 3360 -692 5924 -685
rect 3362 -701 3428 -692
rect 962 -944 992 -918
rect 1162 -944 1192 -918
rect 1364 -944 1394 -918
rect 1564 -944 1594 -918
rect 3380 -732 3410 -701
rect 3476 -732 3506 -692
rect 3554 -701 3620 -692
rect 3572 -732 3602 -701
rect 3668 -732 3698 -692
rect 3746 -701 3812 -692
rect 3764 -732 3794 -701
rect 3860 -732 3890 -692
rect 3938 -701 4004 -692
rect 3956 -732 3986 -701
rect 4052 -732 4082 -692
rect 4130 -701 4196 -692
rect 4148 -732 4178 -701
rect 4244 -732 4274 -692
rect 4322 -701 4388 -692
rect 4340 -732 4370 -701
rect 4436 -732 4466 -692
rect 4514 -701 4580 -692
rect 4532 -732 4562 -701
rect 4628 -732 4658 -692
rect 4706 -701 4772 -692
rect 4724 -732 4754 -701
rect 4820 -732 4850 -692
rect 4898 -701 4964 -692
rect 4916 -732 4946 -701
rect 5012 -732 5042 -692
rect 5090 -701 5156 -692
rect 5108 -732 5138 -701
rect 5204 -732 5234 -692
rect 5282 -701 5348 -692
rect 5300 -732 5330 -701
rect 5396 -732 5426 -692
rect 5474 -701 5540 -692
rect 5492 -732 5522 -701
rect 5588 -732 5618 -692
rect 5666 -701 5732 -692
rect 5684 -732 5714 -701
rect 5780 -732 5810 -692
rect 5858 -701 5924 -692
rect 5876 -732 5906 -701
rect 594 -996 788 -986
rect 594 -1034 610 -996
rect 772 -1034 788 -996
rect 594 -1046 788 -1034
rect 1994 -1008 2024 -962
rect 2090 -993 2120 -962
rect 2072 -1008 2138 -993
rect 2186 -1008 2216 -962
rect 1994 -1009 2216 -1008
rect 1994 -1043 2088 -1009
rect 2122 -1043 2216 -1009
rect 1994 -1044 2216 -1043
rect 2402 -1010 2432 -962
rect 2498 -993 2528 -962
rect 2480 -1009 2546 -993
rect 2480 -1010 2496 -1009
rect 2402 -1043 2496 -1010
rect 2530 -1010 2546 -1009
rect 2594 -1010 2624 -962
rect 2690 -993 2720 -962
rect 2672 -1009 2738 -993
rect 2672 -1010 2688 -1009
rect 2530 -1043 2688 -1010
rect 2722 -1010 2738 -1009
rect 2786 -1010 2816 -962
rect 2882 -993 2912 -962
rect 2864 -1009 2930 -993
rect 2864 -1010 2880 -1009
rect 2722 -1043 2880 -1010
rect 2914 -1010 2930 -1009
rect 2978 -1010 3008 -962
rect 3074 -993 3104 -962
rect 3056 -1009 3122 -993
rect 3056 -1010 3072 -1009
rect 2914 -1043 3072 -1010
rect 3106 -1010 3122 -1009
rect 3170 -1010 3200 -962
rect 3106 -1043 3200 -1010
rect 3380 -1042 3410 -984
rect 3476 -1015 3506 -984
rect 3458 -1031 3524 -1015
rect 3458 -1042 3474 -1031
rect 2402 -1044 3200 -1043
rect 2072 -1059 2138 -1044
rect 2480 -1059 2546 -1044
rect 2672 -1059 2738 -1044
rect 2864 -1059 2930 -1044
rect 3056 -1059 3122 -1044
rect 3378 -1065 3474 -1042
rect 3508 -1042 3524 -1031
rect 3572 -1042 3602 -984
rect 3668 -1015 3698 -984
rect 3650 -1031 3716 -1015
rect 3650 -1042 3666 -1031
rect 3508 -1065 3666 -1042
rect 3700 -1042 3716 -1031
rect 3764 -1042 3794 -984
rect 3860 -1015 3890 -984
rect 3842 -1031 3908 -1015
rect 3842 -1042 3858 -1031
rect 3700 -1065 3858 -1042
rect 3892 -1042 3908 -1031
rect 3956 -1042 3986 -984
rect 4052 -1015 4082 -984
rect 4034 -1031 4100 -1015
rect 4034 -1042 4050 -1031
rect 3892 -1065 4050 -1042
rect 4084 -1042 4100 -1031
rect 4148 -1042 4178 -984
rect 4244 -1015 4274 -984
rect 4226 -1031 4292 -1015
rect 4226 -1042 4242 -1031
rect 4084 -1065 4242 -1042
rect 4276 -1042 4292 -1031
rect 4340 -1042 4370 -984
rect 4436 -1015 4466 -984
rect 4418 -1031 4484 -1015
rect 4418 -1042 4434 -1031
rect 4276 -1065 4434 -1042
rect 4468 -1042 4484 -1031
rect 4532 -1042 4562 -984
rect 4628 -1015 4658 -984
rect 4610 -1031 4676 -1015
rect 4610 -1042 4626 -1031
rect 4468 -1065 4626 -1042
rect 4660 -1042 4676 -1031
rect 4724 -1042 4754 -984
rect 4820 -1015 4850 -984
rect 4802 -1031 4868 -1015
rect 4802 -1042 4818 -1031
rect 4660 -1065 4818 -1042
rect 4852 -1042 4868 -1031
rect 4916 -1042 4946 -984
rect 5012 -1015 5042 -984
rect 4994 -1031 5060 -1015
rect 4994 -1042 5010 -1031
rect 4852 -1065 5010 -1042
rect 5044 -1042 5060 -1031
rect 5108 -1042 5138 -984
rect 5204 -1015 5234 -984
rect 5186 -1031 5252 -1015
rect 5186 -1042 5202 -1031
rect 5044 -1065 5202 -1042
rect 5236 -1042 5252 -1031
rect 5300 -1042 5330 -984
rect 5396 -1015 5426 -984
rect 5378 -1031 5444 -1015
rect 5378 -1042 5394 -1031
rect 5236 -1065 5394 -1042
rect 5428 -1042 5444 -1031
rect 5492 -1042 5522 -984
rect 5588 -1015 5618 -984
rect 5570 -1031 5636 -1015
rect 5570 -1042 5586 -1031
rect 5428 -1065 5586 -1042
rect 5620 -1042 5636 -1031
rect 5684 -1042 5714 -984
rect 5780 -1015 5810 -984
rect 5762 -1031 5828 -1015
rect 5762 -1042 5778 -1031
rect 5620 -1065 5778 -1042
rect 5812 -1042 5828 -1031
rect 5876 -1042 5906 -984
rect 5812 -1065 5908 -1042
rect 3378 -1074 5908 -1065
rect 3458 -1081 3524 -1074
rect 3650 -1081 3716 -1074
rect 3842 -1081 3908 -1074
rect 4034 -1081 4100 -1074
rect 4226 -1081 4292 -1074
rect 4418 -1081 4484 -1074
rect 4610 -1081 4676 -1074
rect 4724 -1078 4754 -1074
rect 4802 -1081 4868 -1074
rect 4994 -1081 5060 -1074
rect 5186 -1081 5252 -1074
rect 5378 -1081 5444 -1074
rect 5570 -1081 5636 -1074
rect 5762 -1081 5828 -1074
<< polycont >>
rect 638 604 778 638
rect -28 136 72 180
rect 146 140 272 180
rect 440 140 570 180
rect 848 144 946 206
rect 1046 138 1144 212
rect 1246 140 1344 214
rect 1446 140 1544 214
rect 1664 138 1926 176
rect 2298 148 2370 190
rect 3264 130 3384 166
rect 354 -122 770 -86
rect 360 -302 780 -248
rect 1988 -360 2022 -326
rect 2180 -360 2214 -326
rect -40 -576 272 -534
rect 432 -576 570 -534
rect 2402 -360 2436 -326
rect 2594 -360 2628 -326
rect 2786 -360 2820 -326
rect 2978 -360 3012 -326
rect 3170 -360 3204 -326
rect 3378 -360 3412 -326
rect 3570 -360 3604 -326
rect 3762 -360 3796 -326
rect 3954 -360 3988 -326
rect 4146 -360 4180 -326
rect 4338 -360 4372 -326
rect 4530 -360 4564 -326
rect 4722 -360 4756 -326
rect 4914 -360 4948 -326
rect 5106 -360 5140 -326
rect 5298 -360 5332 -326
rect 5490 -360 5524 -326
rect 5682 -360 5716 -326
rect 5874 -360 5908 -326
rect 844 -568 948 -530
rect 1052 -610 1150 -536
rect 1252 -612 1350 -538
rect 1452 -612 1550 -538
rect 1698 -576 1858 -518
rect 2084 -554 2118 -520
rect 2296 -582 2392 -548
rect 2498 -554 2532 -520
rect 2690 -554 2724 -520
rect 2882 -554 2916 -520
rect 3074 -554 3108 -520
rect 3270 -570 3374 -532
rect 3474 -554 3508 -520
rect 3666 -554 3700 -520
rect 3858 -554 3892 -520
rect 4050 -554 4084 -520
rect 4242 -554 4276 -520
rect 4434 -554 4468 -520
rect 4626 -554 4660 -520
rect 4818 -554 4852 -520
rect 5010 -554 5044 -520
rect 5202 -554 5236 -520
rect 5394 -554 5428 -520
rect 5586 -554 5620 -520
rect 5778 -554 5812 -520
rect 1992 -663 2026 -629
rect 2184 -663 2218 -629
rect 2400 -663 2434 -629
rect 2592 -663 2626 -629
rect 2784 -663 2818 -629
rect 2976 -663 3010 -629
rect 3168 -663 3202 -629
rect 3378 -685 3412 -651
rect 3570 -685 3604 -651
rect 3762 -685 3796 -651
rect 3954 -685 3988 -651
rect 4146 -685 4180 -651
rect 4338 -685 4372 -651
rect 4530 -685 4564 -651
rect 4722 -685 4756 -651
rect 4914 -685 4948 -651
rect 5106 -685 5140 -651
rect 5298 -685 5332 -651
rect 5490 -685 5524 -651
rect 5682 -685 5716 -651
rect 5874 -685 5908 -651
rect 610 -1034 772 -996
rect 2088 -1043 2122 -1009
rect 2496 -1043 2530 -1009
rect 2688 -1043 2722 -1009
rect 2880 -1043 2914 -1009
rect 3072 -1043 3106 -1009
rect 3474 -1065 3508 -1031
rect 3666 -1065 3700 -1031
rect 3858 -1065 3892 -1031
rect 4050 -1065 4084 -1031
rect 4242 -1065 4276 -1031
rect 4434 -1065 4468 -1031
rect 4626 -1065 4660 -1031
rect 4818 -1065 4852 -1031
rect 5010 -1065 5044 -1031
rect 5202 -1065 5236 -1031
rect 5394 -1065 5428 -1031
rect 5586 -1065 5620 -1031
rect 5778 -1065 5812 -1031
<< locali >>
rect 2228 658 2322 670
rect 618 646 792 654
rect 618 638 794 646
rect 618 604 638 638
rect 778 604 794 638
rect 2228 624 2240 658
rect 2308 650 2322 658
rect 2308 624 2548 650
rect 2228 616 2548 624
rect 2232 614 2320 616
rect -152 578 -86 596
rect 618 592 794 604
rect 618 588 792 592
rect -152 290 -138 578
rect -100 290 -86 578
rect 510 506 544 522
rect -152 272 -86 290
rect 298 272 332 332
rect 298 238 428 272
rect 510 262 544 278
rect 598 506 632 522
rect 598 262 632 278
rect 710 506 744 522
rect 798 520 832 522
rect 794 506 832 520
rect 794 278 798 506
rect 710 262 744 278
rect 794 266 832 278
rect 798 262 832 266
rect -136 180 88 198
rect 72 136 88 180
rect -136 122 88 136
rect 134 180 286 200
rect 134 140 146 180
rect 272 140 286 180
rect 134 122 286 140
rect 386 198 428 238
rect 832 206 964 220
rect 386 180 586 198
rect 386 140 440 180
rect 570 140 586 180
rect -136 120 86 122
rect 386 120 586 140
rect 832 144 848 206
rect 946 144 964 206
rect 832 132 964 144
rect 1030 212 1160 226
rect 1030 138 1046 212
rect 1144 138 1160 212
rect 1030 124 1160 138
rect 1222 214 1362 230
rect 1222 140 1246 214
rect 1344 140 1362 214
rect 1222 122 1362 140
rect 1428 214 1564 230
rect 1428 140 1446 214
rect 1544 140 1564 214
rect 1428 122 1564 140
rect 1648 176 1946 192
rect 1648 138 1664 176
rect 1926 138 1946 176
rect 2272 190 2386 198
rect 2272 148 2298 190
rect 2370 148 2386 190
rect 2272 140 2386 148
rect 3246 166 3400 182
rect 1648 126 1946 138
rect 3246 130 3264 166
rect 3384 130 3400 166
rect 3246 124 3400 130
rect 386 80 428 120
rect 386 12 420 80
rect 510 70 544 86
rect 510 -6 544 10
rect 598 70 632 86
rect 598 -6 632 10
rect 710 70 744 86
rect 710 -6 744 10
rect 798 70 832 86
rect 798 -6 832 10
rect 338 -86 792 -74
rect 338 -122 354 -86
rect 770 -122 792 -86
rect 338 -132 792 -122
rect 344 -248 798 -236
rect 344 -302 360 -248
rect 780 -302 798 -248
rect 344 -312 798 -302
rect 3362 -326 5924 -324
rect 1972 -360 1988 -326
rect 2022 -360 2038 -326
rect 2164 -360 2180 -326
rect 2214 -360 2230 -326
rect 2386 -360 2402 -326
rect 2436 -360 2452 -326
rect 2578 -360 2594 -326
rect 2628 -360 2644 -326
rect 2770 -360 2786 -326
rect 2820 -360 2836 -326
rect 2962 -360 2978 -326
rect 3012 -360 3028 -326
rect 3154 -360 3170 -326
rect 3204 -360 3220 -326
rect 3362 -360 3378 -326
rect 3412 -360 3570 -326
rect 3604 -360 3762 -326
rect 3796 -360 3954 -326
rect 3988 -360 4146 -326
rect 4180 -360 4338 -326
rect 4372 -360 4530 -326
rect 4564 -360 4722 -326
rect 4756 -360 4914 -326
rect 4948 -360 5106 -326
rect 5140 -360 5298 -326
rect 5332 -360 5490 -326
rect 5524 -360 5682 -326
rect 5716 -360 5874 -326
rect 5908 -360 5924 -326
rect 32 -412 102 -388
rect 32 -460 48 -412
rect 86 -460 102 -412
rect 32 -486 102 -460
rect 210 -406 244 -390
rect 210 -482 244 -466
rect 298 -406 332 -390
rect 298 -482 332 -466
rect 386 -406 420 -390
rect 386 -514 420 -466
rect 510 -404 544 -388
rect 510 -480 544 -464
rect 598 -404 632 -388
rect 598 -480 632 -464
rect 710 -404 744 -388
rect 710 -480 744 -464
rect 798 -404 832 -388
rect 798 -480 832 -464
rect 916 -408 950 -392
rect 916 -484 950 -468
rect 1004 -408 1038 -392
rect 1004 -484 1038 -468
rect 1116 -410 1150 -394
rect 1116 -486 1150 -470
rect 1204 -410 1238 -394
rect 1204 -486 1238 -470
rect 1318 -408 1352 -392
rect 1318 -484 1352 -468
rect 1406 -408 1440 -392
rect 1406 -484 1440 -468
rect 1518 -410 1552 -394
rect 1518 -486 1552 -470
rect 1606 -410 1640 -394
rect 1606 -486 1640 -470
rect 1940 -410 1974 -394
rect 1940 -486 1974 -470
rect 2036 -410 2070 -394
rect 2036 -486 2070 -470
rect 2132 -410 2166 -394
rect 2132 -486 2166 -470
rect 2228 -410 2262 -394
rect 2228 -486 2262 -470
rect 2354 -410 2388 -394
rect 2354 -486 2388 -470
rect 2450 -410 2484 -394
rect 2450 -486 2484 -470
rect 2546 -410 2580 -394
rect 2546 -486 2580 -470
rect 2642 -410 2676 -394
rect 2642 -486 2676 -470
rect 2738 -410 2772 -394
rect 2738 -486 2772 -470
rect 2834 -410 2868 -394
rect 2834 -486 2868 -470
rect 2930 -410 2964 -394
rect 2930 -486 2964 -470
rect 3026 -410 3060 -394
rect 3026 -486 3060 -470
rect 3122 -410 3156 -394
rect 3122 -486 3156 -470
rect 3218 -410 3252 -394
rect 3218 -486 3252 -470
rect 3330 -410 3364 -394
rect 3330 -486 3364 -470
rect 3426 -410 3460 -394
rect 3426 -486 3460 -470
rect 3522 -410 3556 -394
rect 3522 -486 3556 -470
rect 3618 -410 3652 -394
rect 3618 -486 3652 -470
rect 3714 -410 3748 -394
rect 3714 -486 3748 -470
rect 3810 -410 3844 -394
rect 3810 -486 3844 -470
rect 3906 -410 3940 -394
rect 3906 -486 3940 -470
rect 4002 -410 4036 -394
rect 4002 -486 4036 -470
rect 4098 -410 4132 -394
rect 4098 -486 4132 -470
rect 4194 -410 4228 -394
rect 4194 -486 4228 -470
rect 4290 -410 4324 -394
rect 4290 -486 4324 -470
rect 4386 -410 4420 -394
rect 4386 -486 4420 -470
rect 4482 -410 4516 -394
rect 4482 -486 4516 -470
rect 4578 -410 4612 -394
rect 4578 -486 4612 -470
rect 4674 -410 4708 -394
rect 4674 -486 4708 -470
rect 4770 -410 4804 -394
rect 4770 -486 4804 -470
rect 4866 -410 4900 -394
rect 4866 -486 4900 -470
rect 4962 -410 4996 -394
rect 4962 -486 4996 -470
rect 5058 -410 5092 -394
rect 5058 -486 5092 -470
rect 5154 -410 5188 -394
rect 5154 -486 5188 -470
rect 5250 -410 5284 -394
rect 5250 -486 5284 -470
rect 5346 -410 5380 -394
rect 5346 -486 5380 -470
rect 5442 -410 5476 -394
rect 5442 -486 5476 -470
rect 5538 -410 5572 -394
rect 5538 -486 5572 -470
rect 5634 -410 5668 -394
rect 5634 -486 5668 -470
rect 5730 -410 5764 -394
rect 5730 -486 5764 -470
rect 5826 -410 5860 -394
rect 5826 -486 5860 -470
rect 5922 -410 5956 -394
rect 5922 -486 5956 -470
rect -56 -520 -10 -516
rect 210 -520 286 -516
rect -56 -534 286 -520
rect -56 -576 -40 -534
rect 272 -576 286 -534
rect -56 -592 286 -576
rect 210 -594 286 -592
rect 386 -534 586 -514
rect 1678 -518 1876 -506
rect 386 -576 432 -534
rect 570 -576 586 -534
rect 386 -594 586 -576
rect 828 -530 968 -518
rect 828 -568 844 -530
rect 948 -568 968 -530
rect 828 -580 968 -568
rect 1036 -536 1166 -522
rect 386 -632 420 -594
rect 1036 -610 1052 -536
rect 1150 -610 1166 -536
rect 1036 -624 1166 -610
rect 1228 -538 1368 -520
rect 1228 -612 1252 -538
rect 1350 -612 1368 -538
rect 1228 -628 1368 -612
rect 1434 -538 1570 -520
rect 1434 -612 1452 -538
rect 1550 -612 1570 -538
rect 1678 -576 1698 -518
rect 1858 -576 1876 -518
rect 2068 -554 2084 -520
rect 2118 -554 2134 -520
rect 2268 -548 2424 -542
rect 1678 -588 1876 -576
rect 2268 -582 2296 -548
rect 2392 -582 2424 -548
rect 2482 -554 2498 -520
rect 2532 -554 2548 -520
rect 2674 -554 2690 -520
rect 2724 -554 2740 -520
rect 2866 -554 2882 -520
rect 2916 -554 2932 -520
rect 3058 -554 3074 -520
rect 3108 -554 3124 -520
rect 3252 -532 3474 -520
rect 3252 -570 3270 -532
rect 3374 -554 3474 -532
rect 3508 -554 3666 -520
rect 3700 -554 3858 -520
rect 3892 -554 4050 -520
rect 4084 -554 4242 -520
rect 4276 -554 4434 -520
rect 4468 -554 4626 -520
rect 4660 -554 4818 -520
rect 4852 -554 5010 -520
rect 5044 -554 5202 -520
rect 5236 -554 5394 -520
rect 5428 -554 5586 -520
rect 5620 -554 5778 -520
rect 5812 -554 5908 -520
rect 3374 -556 5908 -554
rect 3374 -570 3400 -556
rect 3252 -582 3400 -570
rect 2268 -594 2424 -582
rect 1434 -628 1570 -612
rect 298 -666 420 -632
rect 6 -732 72 -716
rect 6 -928 22 -732
rect 56 -928 72 -732
rect 6 -946 72 -928
rect 210 -720 244 -704
rect 210 -964 244 -948
rect 298 -720 332 -666
rect 510 -672 544 -656
rect 298 -964 332 -948
rect 386 -720 420 -702
rect 510 -916 544 -900
rect 598 -672 632 -656
rect 598 -916 632 -900
rect 710 -672 744 -656
rect 710 -916 744 -900
rect 798 -672 832 -656
rect 798 -916 832 -900
rect 916 -678 950 -662
rect 916 -922 950 -906
rect 1004 -678 1038 -662
rect 1004 -922 1038 -906
rect 1116 -678 1150 -662
rect 1116 -922 1150 -906
rect 1204 -678 1238 -662
rect 1204 -922 1238 -906
rect 1318 -678 1352 -662
rect 1318 -922 1352 -906
rect 1406 -678 1440 -662
rect 1406 -922 1440 -906
rect 1518 -678 1552 -662
rect 1518 -922 1552 -906
rect 1606 -678 1640 -662
rect 1976 -663 1992 -629
rect 2026 -663 2042 -629
rect 2168 -663 2184 -629
rect 2218 -663 2234 -629
rect 2384 -663 2400 -629
rect 2434 -663 2450 -629
rect 2576 -663 2592 -629
rect 2626 -663 2642 -629
rect 2768 -663 2784 -629
rect 2818 -663 2834 -629
rect 2960 -663 2976 -629
rect 3010 -663 3026 -629
rect 3152 -663 3168 -629
rect 3202 -663 3218 -629
rect 5872 -651 5908 -556
rect 3362 -685 3378 -651
rect 3412 -658 3428 -651
rect 3554 -658 3570 -651
rect 3412 -685 3570 -658
rect 3604 -658 3620 -651
rect 3746 -658 3762 -651
rect 3604 -685 3762 -658
rect 3796 -658 3812 -651
rect 3938 -658 3954 -651
rect 3796 -685 3954 -658
rect 3988 -658 4004 -651
rect 4130 -658 4146 -651
rect 3988 -685 4146 -658
rect 4180 -658 4196 -651
rect 4322 -658 4338 -651
rect 4180 -685 4338 -658
rect 4372 -658 4388 -651
rect 4514 -658 4530 -651
rect 4372 -685 4530 -658
rect 4564 -658 4580 -651
rect 4706 -658 4722 -651
rect 4564 -685 4722 -658
rect 4756 -658 4772 -651
rect 4898 -658 4914 -651
rect 4756 -685 4914 -658
rect 4948 -658 4964 -651
rect 5090 -658 5106 -651
rect 4948 -685 5106 -658
rect 5140 -658 5156 -651
rect 5282 -658 5298 -651
rect 5140 -685 5298 -658
rect 5332 -658 5348 -651
rect 5474 -658 5490 -651
rect 5332 -685 5490 -658
rect 5524 -658 5540 -651
rect 5666 -658 5682 -651
rect 5524 -685 5682 -658
rect 5716 -658 5732 -651
rect 5858 -658 5874 -651
rect 5716 -685 5874 -658
rect 5908 -685 5924 -651
rect 3362 -694 5908 -685
rect 1606 -922 1640 -906
rect 1944 -722 1978 -706
rect 386 -964 420 -948
rect 1944 -966 1978 -950
rect 2040 -722 2074 -706
rect 2040 -966 2074 -950
rect 2136 -722 2170 -706
rect 2136 -966 2170 -950
rect 2232 -722 2266 -706
rect 2232 -966 2266 -950
rect 2352 -722 2386 -706
rect 2352 -966 2386 -950
rect 2448 -722 2482 -706
rect 2448 -966 2482 -950
rect 2544 -722 2578 -706
rect 2544 -966 2578 -950
rect 2640 -722 2674 -706
rect 2640 -966 2674 -950
rect 2736 -722 2770 -706
rect 2736 -966 2770 -950
rect 2832 -722 2866 -706
rect 2832 -966 2866 -950
rect 2928 -722 2962 -706
rect 2928 -966 2962 -950
rect 3024 -722 3058 -706
rect 3024 -966 3058 -950
rect 3120 -722 3154 -706
rect 3120 -966 3154 -950
rect 3216 -722 3250 -706
rect 3216 -966 3250 -950
rect 3330 -744 3364 -728
rect 594 -996 788 -986
rect 3330 -988 3364 -972
rect 3426 -744 3460 -728
rect 3426 -988 3460 -972
rect 3522 -744 3556 -728
rect 3522 -988 3556 -972
rect 3618 -744 3652 -728
rect 3618 -988 3652 -972
rect 3714 -744 3748 -728
rect 3714 -988 3748 -972
rect 3810 -744 3844 -728
rect 3810 -988 3844 -972
rect 3906 -744 3940 -728
rect 3906 -988 3940 -972
rect 4002 -744 4036 -728
rect 4002 -988 4036 -972
rect 4098 -744 4132 -728
rect 4098 -988 4132 -972
rect 4194 -744 4228 -728
rect 4194 -988 4228 -972
rect 4290 -744 4324 -728
rect 4290 -988 4324 -972
rect 4386 -744 4420 -728
rect 4386 -988 4420 -972
rect 4482 -744 4516 -728
rect 4482 -988 4516 -972
rect 4578 -744 4612 -728
rect 4578 -988 4612 -972
rect 4674 -744 4708 -728
rect 4674 -988 4708 -972
rect 4770 -744 4804 -728
rect 4770 -988 4804 -972
rect 4866 -744 4900 -728
rect 4866 -988 4900 -972
rect 4962 -744 4996 -728
rect 4962 -988 4996 -972
rect 5058 -744 5092 -728
rect 5058 -988 5092 -972
rect 5154 -744 5188 -728
rect 5154 -988 5188 -972
rect 5250 -744 5284 -728
rect 5250 -988 5284 -972
rect 5346 -744 5380 -728
rect 5346 -988 5380 -972
rect 5442 -744 5476 -728
rect 5442 -988 5476 -972
rect 5538 -744 5572 -728
rect 5538 -988 5572 -972
rect 5634 -744 5668 -728
rect 5634 -988 5668 -972
rect 5730 -744 5764 -728
rect 5730 -988 5764 -972
rect 5826 -744 5860 -728
rect 5826 -988 5860 -972
rect 5922 -744 5956 -728
rect 5922 -988 5956 -972
rect 594 -1034 610 -996
rect 772 -1034 788 -996
rect 594 -1046 788 -1034
rect 2072 -1043 2088 -1009
rect 2122 -1043 2138 -1009
rect 2232 -1012 2320 -1010
rect 2480 -1012 2496 -1009
rect 2228 -1020 2496 -1012
rect 2228 -1054 2240 -1020
rect 2308 -1043 2496 -1020
rect 2530 -1012 2546 -1009
rect 2530 -1043 2548 -1012
rect 2672 -1043 2688 -1009
rect 2722 -1043 2738 -1009
rect 2864 -1043 2880 -1009
rect 2914 -1043 2930 -1009
rect 3056 -1043 3072 -1009
rect 3106 -1043 3122 -1009
rect 3458 -1038 3474 -1031
rect 2308 -1046 2548 -1043
rect 2308 -1054 2322 -1046
rect 2228 -1066 2322 -1054
rect 3378 -1065 3474 -1038
rect 3508 -1040 3524 -1031
rect 3650 -1040 3666 -1031
rect 3508 -1065 3666 -1040
rect 3700 -1040 3716 -1031
rect 3842 -1040 3858 -1031
rect 3700 -1065 3858 -1040
rect 3892 -1040 3908 -1031
rect 4034 -1040 4050 -1031
rect 3892 -1065 4050 -1040
rect 4084 -1040 4100 -1031
rect 4226 -1040 4242 -1031
rect 4084 -1065 4242 -1040
rect 4276 -1040 4292 -1031
rect 4418 -1040 4434 -1031
rect 4276 -1065 4434 -1040
rect 4468 -1040 4484 -1031
rect 4610 -1040 4626 -1031
rect 4468 -1065 4626 -1040
rect 4660 -1040 4676 -1031
rect 4802 -1040 4818 -1031
rect 4660 -1065 4818 -1040
rect 4852 -1040 4868 -1031
rect 4994 -1040 5010 -1031
rect 4852 -1065 5010 -1040
rect 5044 -1040 5060 -1031
rect 5186 -1040 5202 -1031
rect 5044 -1065 5202 -1040
rect 5236 -1040 5252 -1031
rect 5378 -1040 5394 -1031
rect 5236 -1065 5394 -1040
rect 5428 -1040 5444 -1031
rect 5570 -1040 5586 -1031
rect 5428 -1065 5586 -1040
rect 5620 -1040 5636 -1031
rect 5762 -1038 5778 -1031
rect 5746 -1040 5778 -1038
rect 5620 -1065 5778 -1040
rect 5812 -1040 5828 -1031
rect 5812 -1065 5908 -1040
rect 3378 -1072 5908 -1065
rect 3457 -1074 5908 -1072
<< viali >>
rect 638 604 778 638
rect 2240 624 2308 658
rect -138 290 -100 578
rect 510 278 544 506
rect 598 278 632 506
rect 710 278 744 506
rect 744 278 746 506
rect 798 278 832 506
rect -170 136 -28 180
rect -28 136 28 180
rect 146 140 272 180
rect 848 144 946 206
rect 1046 138 1144 212
rect 1246 140 1344 214
rect 1446 140 1544 214
rect 1664 138 1926 176
rect 2298 148 2370 190
rect 3264 130 3384 166
rect 510 10 544 70
rect 598 10 632 70
rect 710 10 744 70
rect 798 10 832 70
rect 354 -122 770 -86
rect 360 -302 780 -248
rect 48 -460 86 -412
rect 210 -466 244 -406
rect 298 -466 332 -406
rect 386 -466 420 -406
rect 510 -464 544 -404
rect 598 -464 632 -404
rect 710 -464 744 -404
rect 798 -464 832 -404
rect 916 -468 950 -408
rect 1004 -468 1038 -408
rect 1116 -470 1150 -410
rect 1204 -470 1238 -410
rect 1318 -468 1352 -408
rect 1406 -468 1440 -408
rect 1518 -470 1552 -410
rect 1606 -470 1640 -410
rect 1940 -470 1974 -410
rect 2036 -470 2070 -410
rect 2132 -470 2166 -410
rect 2228 -470 2262 -410
rect 2354 -470 2388 -410
rect 2450 -470 2484 -410
rect 2546 -470 2580 -410
rect 2642 -470 2676 -410
rect 2738 -470 2772 -410
rect 2834 -470 2868 -410
rect 2930 -470 2964 -410
rect 3026 -470 3060 -410
rect 3122 -470 3156 -410
rect 3218 -470 3252 -410
rect 3330 -470 3364 -410
rect 3426 -470 3460 -410
rect 3522 -470 3556 -410
rect 3618 -470 3652 -410
rect 3714 -470 3748 -410
rect 3810 -470 3844 -410
rect 3906 -470 3940 -410
rect 4002 -470 4036 -410
rect 4098 -470 4132 -410
rect 4194 -470 4228 -410
rect 4290 -470 4324 -410
rect 4386 -470 4420 -410
rect 4482 -470 4516 -410
rect 4578 -470 4612 -410
rect 4674 -470 4708 -410
rect 4770 -470 4804 -410
rect 4866 -470 4900 -410
rect 4962 -470 4996 -410
rect 5058 -470 5092 -410
rect 5154 -470 5188 -410
rect 5250 -470 5284 -410
rect 5346 -470 5380 -410
rect 5442 -470 5476 -410
rect 5538 -470 5572 -410
rect 5634 -470 5668 -410
rect 5730 -470 5764 -410
rect 5826 -470 5860 -410
rect 5922 -470 5956 -410
rect -40 -576 272 -534
rect 844 -568 948 -530
rect 1052 -610 1150 -536
rect 1252 -612 1350 -538
rect 1452 -612 1550 -538
rect 1698 -576 1858 -518
rect 2296 -582 2392 -548
rect 3270 -570 3374 -532
rect 22 -928 56 -732
rect 210 -948 244 -720
rect 298 -948 332 -720
rect 386 -948 420 -720
rect 510 -900 544 -672
rect 598 -900 632 -672
rect 710 -900 744 -672
rect 798 -900 832 -672
rect 916 -906 950 -678
rect 1004 -906 1038 -678
rect 1116 -906 1150 -678
rect 1204 -906 1238 -678
rect 1318 -906 1352 -678
rect 1406 -906 1440 -678
rect 1518 -906 1552 -678
rect 1606 -906 1640 -678
rect 1944 -950 1978 -722
rect 2040 -950 2074 -722
rect 2136 -950 2170 -722
rect 2232 -950 2266 -722
rect 2352 -950 2386 -722
rect 2448 -950 2482 -722
rect 2544 -950 2578 -722
rect 2640 -950 2674 -722
rect 2736 -950 2770 -722
rect 2832 -950 2866 -722
rect 2928 -950 2962 -722
rect 3024 -950 3058 -722
rect 3120 -950 3154 -722
rect 3216 -950 3250 -722
rect 3330 -972 3364 -744
rect 3426 -972 3460 -744
rect 3522 -972 3556 -744
rect 3618 -972 3652 -744
rect 3714 -972 3748 -744
rect 3810 -972 3844 -744
rect 3906 -972 3940 -744
rect 4002 -972 4036 -744
rect 4098 -972 4132 -744
rect 4194 -972 4228 -744
rect 4290 -972 4324 -744
rect 4386 -972 4420 -744
rect 4482 -972 4516 -744
rect 4578 -972 4612 -744
rect 4674 -972 4708 -744
rect 4770 -972 4804 -744
rect 4866 -972 4900 -744
rect 4962 -972 4996 -744
rect 5058 -972 5092 -744
rect 5154 -972 5188 -744
rect 5250 -972 5284 -744
rect 5346 -972 5380 -744
rect 5442 -972 5476 -744
rect 5538 -972 5572 -744
rect 5634 -972 5668 -744
rect 5730 -972 5764 -744
rect 5826 -972 5860 -744
rect 5922 -972 5956 -744
rect 610 -1034 772 -998
rect 2240 -1054 2308 -1020
<< metal1 >>
rect -280 1208 6008 1268
rect -280 766 -188 1208
rect 5906 766 6008 1208
rect -280 698 6008 766
rect -278 -1080 -213 698
rect -152 616 -84 698
rect -152 578 -86 616
rect -152 290 -138 578
rect -100 290 -86 578
rect 12 456 42 698
rect 210 630 242 698
rect 384 636 424 698
rect 212 464 242 630
rect 386 468 422 636
rect 512 634 544 698
rect 600 646 792 654
rect 600 638 794 646
rect 512 518 542 634
rect 600 604 638 638
rect 778 604 794 638
rect 600 592 794 604
rect 600 588 792 592
rect 600 550 632 588
rect 1930 568 1980 698
rect 2228 658 2322 670
rect 2228 624 2240 658
rect 2308 624 2322 658
rect 2228 616 2322 624
rect 2232 614 2320 616
rect 598 518 632 550
rect 1924 556 2002 568
rect 488 508 564 518
rect -152 272 -86 290
rect 488 276 502 508
rect 558 276 564 508
rect 98 202 132 274
rect 488 266 564 276
rect 592 506 638 518
rect 592 278 598 506
rect 632 278 638 506
rect 592 266 638 278
rect 696 506 756 518
rect 98 198 256 202
rect -182 186 40 198
rect -182 132 -170 186
rect 28 132 40 186
rect -182 120 40 132
rect 98 180 286 198
rect 98 140 146 180
rect 272 140 286 180
rect 98 120 286 140
rect -137 119 9 120
rect -137 118 -59 119
rect 98 118 132 120
rect -2 70 56 82
rect -2 10 0 70
rect 54 10 56 70
rect 98 56 130 118
rect 598 82 632 266
rect 696 264 756 278
rect 792 506 838 520
rect 792 278 798 506
rect 832 278 838 506
rect 792 266 838 278
rect 890 506 962 522
rect 890 282 900 506
rect 956 282 962 506
rect 998 498 1034 524
rect 1088 508 1160 524
rect 890 266 962 282
rect 798 220 832 266
rect 998 228 1032 290
rect 1088 280 1100 508
rect 1156 280 1160 508
rect 1198 490 1234 524
rect 1290 508 1362 522
rect 1088 268 1160 280
rect 1198 230 1232 292
rect 1290 280 1302 508
rect 1358 280 1362 508
rect 1400 494 1436 524
rect 1490 508 1562 522
rect 1290 266 1362 280
rect 1400 230 1434 288
rect 1490 280 1502 508
rect 1558 280 1562 508
rect 1600 494 1634 524
rect 1924 326 1934 556
rect 1990 326 2002 556
rect 2114 554 2192 566
rect 1924 314 2002 326
rect 1490 266 1562 280
rect 798 216 964 220
rect 796 206 964 216
rect 796 186 848 206
rect 798 144 848 186
rect 946 180 964 206
rect 998 212 1170 228
rect 946 144 966 180
rect 798 132 966 144
rect 998 138 1046 212
rect 1144 138 1170 212
rect 798 82 832 132
rect 998 120 1170 138
rect 1198 214 1362 230
rect 1198 140 1246 214
rect 1344 140 1362 214
rect 1198 122 1362 140
rect 1400 214 1566 230
rect 1400 140 1446 214
rect 1544 140 1566 214
rect 1400 122 1566 140
rect 1600 192 1634 290
rect 2038 238 2074 348
rect 2114 326 2126 554
rect 2180 326 2192 554
rect 2232 538 2266 614
rect 2332 554 2404 566
rect 2114 312 2192 326
rect 2230 242 2266 338
rect 2332 326 2340 554
rect 2396 326 2404 554
rect 2528 554 2600 564
rect 2332 312 2404 326
rect 2036 204 2074 238
rect 2228 204 2266 242
rect 1600 176 1946 192
rect 1600 138 1664 176
rect 1926 138 1946 176
rect 1600 124 1946 138
rect 2036 190 2384 204
rect 2036 168 2298 190
rect 504 80 550 82
rect 200 72 254 80
rect -2 -2 56 10
rect 200 -2 254 12
rect 500 70 554 80
rect 500 -2 554 10
rect 592 70 638 82
rect 704 80 750 82
rect 592 10 598 70
rect 632 10 638 70
rect 592 -2 638 10
rect 700 70 754 80
rect 700 -2 754 10
rect 792 70 838 82
rect 792 10 798 70
rect 832 10 838 70
rect 792 -2 838 10
rect 896 70 958 84
rect 896 10 900 70
rect 952 10 958 70
rect 998 64 1032 120
rect 1096 72 1158 84
rect 896 -2 958 10
rect 1096 12 1100 72
rect 1152 12 1158 72
rect 1198 66 1232 122
rect 1298 70 1360 84
rect 1096 -2 1158 12
rect 1298 10 1304 70
rect 1356 10 1360 70
rect 1400 62 1434 122
rect 1600 112 1636 124
rect 1498 72 1560 84
rect 1298 -2 1360 10
rect 1498 12 1504 72
rect 1556 12 1560 72
rect 1600 64 1634 112
rect 1498 -2 1560 12
rect 338 -78 792 -66
rect 338 -130 354 -78
rect 772 -130 792 -78
rect 338 -132 792 -130
rect 1764 -236 1840 124
rect 1928 74 1990 86
rect 1928 14 1930 74
rect 1986 14 1990 74
rect 2036 64 2072 168
rect 2228 148 2298 168
rect 2370 148 2384 190
rect 2228 138 2384 148
rect 2450 202 2486 342
rect 2528 326 2534 554
rect 2590 326 2600 554
rect 2718 554 2790 566
rect 2528 314 2600 326
rect 2640 202 2676 366
rect 2718 326 2724 554
rect 2780 326 2790 554
rect 2912 552 2984 564
rect 2718 316 2790 326
rect 2830 202 2866 376
rect 2912 324 2918 552
rect 2974 324 2984 552
rect 3100 554 3172 566
rect 2912 314 2984 324
rect 3022 202 3058 406
rect 3100 326 3110 554
rect 3166 326 3172 554
rect 3100 316 3172 326
rect 3210 202 3258 356
rect 2450 182 3258 202
rect 2450 166 3400 182
rect 2118 74 2180 86
rect 1928 0 1990 14
rect 2118 14 2122 74
rect 2178 14 2180 74
rect 2228 54 2264 138
rect 2340 74 2400 86
rect 2118 0 2180 14
rect 2340 14 2344 74
rect 2398 14 2400 74
rect 2450 26 2486 166
rect 2534 74 2594 86
rect 2340 2 2400 14
rect 2534 14 2536 74
rect 2590 14 2594 74
rect 2640 44 2676 166
rect 2726 74 2786 86
rect 2534 2 2594 14
rect 2726 14 2728 74
rect 2782 14 2786 74
rect 2830 34 2866 166
rect 2916 74 2980 86
rect 2726 2 2786 14
rect 2916 14 2920 74
rect 2974 14 2980 74
rect 3024 32 3060 166
rect 3210 130 3264 166
rect 3384 130 3400 166
rect 3210 124 3400 130
rect 3108 74 3172 86
rect 2916 2 2980 14
rect 3108 14 3114 74
rect 3168 14 3172 74
rect 3210 48 3258 124
rect 3108 2 3172 14
rect 3330 -100 3364 34
rect 3521 -100 3555 41
rect 3713 -100 3747 35
rect 3905 -100 3939 35
rect 4099 -100 4133 49
rect 4289 -100 4323 43
rect 4481 -100 4515 51
rect 4673 -100 4707 39
rect 4867 -100 4901 33
rect 5057 -100 5091 33
rect 5251 -100 5285 39
rect 5439 -100 5473 37
rect 5633 -100 5667 31
rect 5827 -100 5861 41
rect 3330 -134 6003 -100
rect 344 -248 1840 -236
rect 344 -302 360 -248
rect 780 -302 1840 -248
rect 344 -312 1840 -302
rect 3318 -276 6002 -240
rect 32 -408 102 -388
rect 504 -394 550 -392
rect 204 -396 250 -394
rect 32 -460 40 -408
rect 96 -460 102 -408
rect 32 -486 102 -460
rect 202 -404 254 -396
rect 202 -480 254 -468
rect 292 -406 338 -394
rect 292 -466 298 -406
rect 332 -466 338 -406
rect 292 -478 338 -466
rect 380 -406 426 -394
rect 380 -466 386 -406
rect 420 -466 426 -406
rect 380 -478 426 -466
rect 502 -404 554 -394
rect 502 -476 554 -464
rect 592 -404 638 -392
rect 592 -464 598 -404
rect 632 -464 638 -404
rect 592 -476 638 -464
rect 698 -404 754 -392
rect 698 -464 702 -404
rect 698 -474 754 -464
rect 792 -404 838 -392
rect 792 -464 798 -404
rect 832 -464 838 -404
rect 700 -476 752 -474
rect 792 -476 838 -464
rect 902 -408 964 -396
rect 902 -468 906 -408
rect 958 -468 964 -408
rect 598 -514 632 -476
rect -54 -516 286 -514
rect -56 -526 286 -516
rect -56 -584 -40 -526
rect 274 -584 286 -526
rect -56 -592 286 -584
rect 598 -592 630 -514
rect 798 -518 832 -476
rect 902 -482 964 -468
rect 998 -408 1044 -396
rect 998 -468 1004 -408
rect 1038 -468 1044 -408
rect 998 -480 1044 -468
rect 1102 -410 1164 -396
rect 1102 -470 1106 -410
rect 1158 -470 1164 -410
rect 1004 -518 1038 -480
rect 1102 -482 1164 -470
rect 1198 -410 1244 -398
rect 1198 -470 1204 -410
rect 1238 -470 1244 -410
rect 1198 -482 1244 -470
rect 1304 -408 1366 -396
rect 1304 -468 1310 -408
rect 1362 -468 1366 -408
rect 1304 -482 1366 -468
rect 1400 -408 1446 -396
rect 1400 -468 1406 -408
rect 1440 -468 1446 -408
rect 1400 -480 1446 -468
rect 1504 -410 1566 -396
rect 1504 -470 1510 -410
rect 1562 -470 1566 -410
rect 798 -530 968 -518
rect 798 -568 844 -530
rect 948 -568 968 -530
rect 798 -580 968 -568
rect 1004 -536 1176 -518
rect 132 -594 210 -592
rect 598 -660 632 -592
rect 798 -660 832 -580
rect 1004 -610 1052 -536
rect 1150 -610 1176 -536
rect 1004 -626 1176 -610
rect 1204 -520 1238 -482
rect 1406 -520 1440 -480
rect 1504 -482 1566 -470
rect 1600 -410 1646 -398
rect 1600 -470 1606 -410
rect 1640 -470 1646 -410
rect 1600 -482 1646 -470
rect 1928 -410 1990 -396
rect 1928 -470 1930 -410
rect 1986 -470 1990 -410
rect 1928 -482 1990 -470
rect 2030 -410 2076 -398
rect 2030 -470 2036 -410
rect 2070 -470 2076 -410
rect 2030 -482 2076 -470
rect 2118 -410 2180 -396
rect 3318 -398 3354 -276
rect 3524 -398 3560 -276
rect 3712 -398 3748 -276
rect 3908 -398 3944 -276
rect 4096 -398 4132 -276
rect 4288 -398 4324 -276
rect 4484 -398 4520 -276
rect 4668 -398 4704 -276
rect 4862 -398 4898 -276
rect 5060 -398 5096 -276
rect 5246 -398 5282 -276
rect 5438 -398 5474 -276
rect 5632 -398 5668 -276
rect 5826 -398 5862 -276
rect 2118 -470 2122 -410
rect 2178 -470 2180 -410
rect 2118 -482 2180 -470
rect 2222 -410 2268 -398
rect 2222 -470 2228 -410
rect 2262 -470 2268 -410
rect 2222 -482 2268 -470
rect 2340 -410 2400 -398
rect 2340 -470 2344 -410
rect 2398 -470 2400 -410
rect 2340 -482 2400 -470
rect 2444 -410 2490 -398
rect 2444 -470 2450 -410
rect 2484 -470 2490 -410
rect 2444 -482 2490 -470
rect 2534 -410 2594 -398
rect 2534 -470 2536 -410
rect 2590 -470 2594 -410
rect 2534 -482 2594 -470
rect 2636 -410 2682 -398
rect 2636 -470 2642 -410
rect 2676 -470 2682 -410
rect 2636 -482 2682 -470
rect 2726 -410 2786 -398
rect 2726 -470 2728 -410
rect 2782 -470 2786 -410
rect 2726 -482 2786 -470
rect 2828 -410 2874 -398
rect 2828 -470 2834 -410
rect 2868 -470 2874 -410
rect 2828 -482 2874 -470
rect 2916 -410 2980 -398
rect 2916 -470 2920 -410
rect 2974 -470 2980 -410
rect 2916 -482 2980 -470
rect 3020 -410 3066 -398
rect 3020 -470 3026 -410
rect 3060 -470 3066 -410
rect 3020 -482 3066 -470
rect 3108 -410 3172 -398
rect 3108 -470 3114 -410
rect 3168 -470 3172 -410
rect 3212 -410 3258 -398
rect 3212 -444 3218 -410
rect 3108 -482 3172 -470
rect 3210 -470 3218 -444
rect 3252 -470 3258 -410
rect 3318 -410 3370 -398
rect 3318 -448 3330 -410
rect 1204 -538 1368 -520
rect 1204 -612 1252 -538
rect 1350 -612 1368 -538
rect 504 -672 550 -660
rect 504 -684 510 -672
rect 490 -696 510 -684
rect 544 -684 550 -672
rect 592 -672 638 -660
rect 544 -696 562 -684
rect 6 -732 72 -716
rect 6 -928 22 -732
rect 56 -928 72 -732
rect 6 -946 72 -928
rect 8 -1080 72 -946
rect 204 -720 250 -708
rect 204 -948 210 -720
rect 244 -948 250 -720
rect 204 -960 250 -948
rect 292 -720 338 -708
rect 292 -948 298 -720
rect 332 -948 338 -720
rect 292 -960 338 -948
rect 380 -720 426 -708
rect 380 -948 386 -720
rect 420 -948 426 -720
rect 490 -900 502 -696
rect 554 -900 562 -696
rect 490 -912 562 -900
rect 592 -900 598 -672
rect 632 -900 638 -672
rect 704 -672 750 -660
rect 704 -684 710 -672
rect 592 -912 638 -900
rect 692 -696 710 -684
rect 744 -684 750 -672
rect 792 -672 838 -660
rect 744 -696 764 -684
rect 692 -900 700 -696
rect 752 -900 764 -696
rect 692 -912 764 -900
rect 792 -900 798 -672
rect 832 -900 838 -672
rect 792 -912 838 -900
rect 896 -678 968 -664
rect 1004 -666 1038 -626
rect 1204 -628 1368 -612
rect 1406 -538 1572 -520
rect 1406 -612 1452 -538
rect 1550 -612 1572 -538
rect 1406 -628 1572 -612
rect 1606 -533 1640 -482
rect 1676 -518 1876 -504
rect 1676 -533 1698 -518
rect 1606 -567 1698 -533
rect 1204 -666 1238 -628
rect 896 -680 916 -678
rect 950 -680 968 -678
rect 896 -904 906 -680
rect 962 -904 968 -680
rect 896 -906 916 -904
rect 950 -906 968 -904
rect 380 -960 426 -948
rect 208 -1080 244 -960
rect 384 -1056 420 -960
rect 382 -1080 420 -1056
rect 510 -1080 546 -912
rect 598 -986 632 -912
rect 708 -914 744 -912
rect 896 -920 968 -906
rect 998 -678 1044 -666
rect 998 -906 1004 -678
rect 1038 -906 1044 -678
rect 998 -918 1044 -906
rect 1094 -678 1166 -666
rect 1094 -906 1106 -678
rect 1162 -906 1166 -678
rect 1004 -922 1040 -918
rect 1094 -922 1166 -906
rect 1198 -678 1244 -666
rect 1198 -906 1204 -678
rect 1238 -906 1244 -678
rect 1198 -918 1244 -906
rect 1296 -678 1368 -664
rect 1406 -666 1440 -628
rect 1296 -906 1308 -678
rect 1364 -906 1368 -678
rect 1204 -922 1240 -918
rect 1296 -920 1368 -906
rect 1400 -678 1446 -666
rect 1400 -906 1406 -678
rect 1440 -906 1446 -678
rect 1400 -918 1446 -906
rect 1496 -678 1568 -664
rect 1606 -666 1640 -567
rect 1676 -576 1698 -567
rect 1858 -533 1876 -518
rect 1858 -567 1989 -533
rect 2036 -564 2072 -482
rect 2228 -540 2264 -482
rect 2228 -548 2404 -540
rect 2228 -564 2296 -548
rect 1858 -576 1876 -567
rect 1676 -586 1876 -576
rect 2036 -582 2296 -564
rect 2392 -582 2404 -548
rect 2036 -592 2404 -582
rect 2450 -561 2484 -482
rect 2641 -561 2675 -482
rect 2831 -561 2865 -482
rect 3029 -561 3063 -482
rect 3210 -520 3258 -470
rect 3324 -470 3330 -448
rect 3364 -470 3370 -410
rect 3324 -482 3370 -470
rect 3416 -410 3474 -398
rect 3472 -470 3474 -410
rect 3416 -484 3474 -470
rect 3516 -410 3562 -398
rect 3516 -470 3522 -410
rect 3556 -470 3562 -410
rect 3516 -482 3562 -470
rect 3608 -410 3666 -398
rect 3664 -470 3666 -410
rect 3608 -484 3666 -470
rect 3708 -410 3754 -398
rect 3708 -470 3714 -410
rect 3748 -470 3754 -410
rect 3708 -482 3754 -470
rect 3798 -410 3856 -398
rect 3854 -470 3856 -410
rect 3798 -484 3856 -470
rect 3900 -410 3946 -398
rect 3900 -470 3906 -410
rect 3940 -470 3946 -410
rect 3900 -482 3946 -470
rect 3990 -410 4048 -398
rect 4046 -470 4048 -410
rect 3990 -484 4048 -470
rect 4092 -410 4138 -398
rect 4092 -470 4098 -410
rect 4132 -470 4138 -410
rect 4092 -482 4138 -470
rect 4180 -410 4238 -398
rect 4180 -470 4182 -410
rect 4180 -484 4238 -470
rect 4284 -410 4330 -398
rect 4284 -470 4290 -410
rect 4324 -470 4330 -410
rect 4284 -482 4330 -470
rect 4374 -410 4432 -398
rect 4430 -470 4432 -410
rect 4374 -484 4432 -470
rect 4476 -410 4522 -398
rect 4476 -470 4482 -410
rect 4516 -470 4522 -410
rect 4476 -482 4522 -470
rect 4566 -410 4624 -398
rect 4622 -470 4624 -410
rect 4566 -484 4624 -470
rect 4668 -410 4714 -398
rect 4668 -470 4674 -410
rect 4708 -470 4714 -410
rect 4668 -482 4714 -470
rect 4760 -410 4818 -398
rect 4816 -470 4818 -410
rect 4760 -484 4818 -470
rect 4860 -410 4906 -398
rect 4860 -470 4866 -410
rect 4900 -470 4906 -410
rect 4860 -482 4906 -470
rect 4952 -410 5010 -398
rect 5008 -470 5010 -410
rect 4952 -484 5010 -470
rect 5052 -410 5098 -398
rect 5052 -470 5058 -410
rect 5092 -470 5098 -410
rect 5052 -482 5098 -470
rect 5142 -410 5200 -398
rect 5198 -470 5200 -410
rect 5142 -484 5200 -470
rect 5244 -410 5290 -398
rect 5244 -470 5250 -410
rect 5284 -470 5290 -410
rect 5244 -482 5290 -470
rect 5336 -410 5394 -398
rect 5392 -470 5394 -410
rect 5336 -484 5394 -470
rect 5436 -410 5482 -398
rect 5436 -470 5442 -410
rect 5476 -470 5482 -410
rect 5436 -482 5482 -470
rect 5526 -410 5584 -398
rect 5582 -470 5584 -410
rect 5526 -484 5584 -470
rect 5628 -410 5674 -398
rect 5628 -470 5634 -410
rect 5668 -470 5674 -410
rect 5628 -482 5674 -470
rect 5718 -410 5776 -398
rect 5774 -470 5776 -410
rect 5718 -484 5776 -470
rect 5820 -410 5866 -398
rect 5820 -470 5826 -410
rect 5860 -470 5866 -410
rect 5820 -482 5866 -470
rect 5910 -410 5968 -398
rect 5966 -470 5968 -410
rect 3210 -532 3394 -520
rect 3210 -561 3270 -532
rect 2450 -570 3270 -561
rect 3374 -570 3394 -532
rect 2450 -582 3394 -570
rect 5826 -556 5862 -482
rect 5910 -484 5968 -470
rect 5922 -486 5956 -484
rect 2036 -600 2266 -592
rect 2036 -634 2074 -600
rect 1496 -906 1508 -678
rect 1564 -906 1568 -678
rect 1406 -922 1442 -918
rect 1496 -920 1568 -906
rect 1600 -678 1646 -666
rect 1600 -906 1606 -678
rect 1640 -906 1646 -678
rect 2038 -710 2074 -634
rect 2228 -638 2266 -600
rect 1600 -918 1646 -906
rect 1924 -722 2002 -710
rect 1606 -922 1640 -918
rect 1924 -952 1934 -722
rect 1990 -952 2002 -722
rect 1924 -964 2002 -952
rect 2034 -722 2080 -710
rect 2034 -950 2040 -722
rect 2074 -950 2080 -722
rect 2034 -962 2080 -950
rect 2114 -722 2192 -708
rect 2230 -710 2266 -638
rect 2450 -595 3258 -582
rect 5826 -592 5964 -556
rect 2114 -950 2126 -722
rect 2180 -950 2192 -722
rect 2114 -962 2192 -950
rect 2226 -722 2272 -710
rect 2226 -950 2232 -722
rect 2266 -950 2272 -722
rect 2226 -962 2272 -950
rect 2332 -722 2404 -708
rect 2450 -710 2484 -595
rect 2643 -710 2677 -595
rect 2825 -710 2859 -595
rect 3025 -710 3059 -595
rect 2332 -950 2340 -722
rect 2396 -950 2404 -722
rect 2332 -962 2404 -950
rect 2442 -722 2488 -710
rect 2442 -950 2448 -722
rect 2482 -950 2488 -722
rect 2442 -962 2488 -950
rect 2528 -722 2600 -710
rect 2528 -950 2534 -722
rect 2590 -950 2600 -722
rect 2528 -960 2600 -950
rect 2634 -722 2680 -710
rect 2730 -712 2776 -710
rect 2634 -950 2640 -722
rect 2674 -950 2680 -722
rect 2538 -962 2584 -960
rect 2634 -962 2680 -950
rect 2718 -722 2790 -712
rect 2718 -950 2724 -722
rect 2780 -950 2790 -722
rect 2825 -722 2872 -710
rect 2825 -785 2832 -722
rect 2718 -962 2790 -950
rect 2826 -950 2832 -785
rect 2866 -950 2872 -722
rect 2826 -962 2872 -950
rect 2912 -720 2984 -710
rect 2912 -948 2918 -720
rect 2974 -948 2984 -720
rect 2912 -950 2928 -948
rect 2962 -950 2984 -948
rect 2912 -960 2984 -950
rect 3018 -722 3064 -710
rect 3114 -712 3160 -710
rect 3018 -950 3024 -722
rect 3058 -950 3064 -722
rect 2922 -962 2968 -960
rect 3018 -962 3064 -950
rect 3100 -722 3172 -712
rect 3100 -950 3110 -722
rect 3166 -950 3172 -722
rect 3100 -962 3172 -950
rect 3210 -722 3258 -595
rect 3210 -950 3216 -722
rect 3250 -752 3258 -722
rect 5928 -724 5964 -592
rect 5922 -732 5964 -724
rect 3324 -744 3370 -732
rect 3420 -740 3466 -732
rect 3250 -950 3256 -752
rect 3210 -962 3256 -950
rect 594 -998 788 -986
rect 594 -1034 610 -998
rect 772 -1034 788 -998
rect 594 -1046 788 -1034
rect -278 -1110 -216 -1080
rect 8 -1110 68 -1080
rect 208 -1110 240 -1080
rect 382 -1110 414 -1080
rect 510 -1110 542 -1080
rect 1934 -1110 1990 -964
rect 2232 -1010 2266 -962
rect 3324 -972 3330 -744
rect 3364 -972 3370 -744
rect 3324 -984 3370 -972
rect 3414 -744 3472 -740
rect 3414 -752 3426 -744
rect 3460 -752 3472 -744
rect 3470 -980 3472 -752
rect 2232 -1012 2320 -1010
rect 2228 -1020 2322 -1012
rect 2228 -1054 2240 -1020
rect 2308 -1054 2322 -1020
rect 2228 -1066 2322 -1054
rect 3330 -1110 3364 -984
rect 3414 -992 3472 -980
rect 3516 -744 3562 -732
rect 3612 -740 3658 -732
rect 3516 -972 3522 -744
rect 3556 -972 3562 -744
rect 3516 -984 3562 -972
rect 3604 -744 3662 -740
rect 3604 -752 3618 -744
rect 3652 -752 3662 -744
rect 3604 -980 3606 -752
rect 3522 -1110 3556 -984
rect 3604 -992 3662 -980
rect 3708 -744 3754 -732
rect 3804 -740 3850 -732
rect 3708 -972 3714 -744
rect 3748 -972 3754 -744
rect 3708 -984 3754 -972
rect 3800 -744 3858 -740
rect 3800 -752 3810 -744
rect 3844 -752 3858 -744
rect 3856 -980 3858 -752
rect 3714 -1110 3748 -984
rect 3800 -992 3858 -980
rect 3900 -744 3946 -732
rect 3996 -740 4042 -732
rect 3900 -972 3906 -744
rect 3940 -972 3946 -744
rect 3900 -984 3946 -972
rect 3992 -744 4050 -740
rect 3992 -752 4002 -744
rect 4036 -752 4050 -744
rect 4048 -980 4050 -752
rect 3906 -1110 3940 -984
rect 3992 -992 4050 -980
rect 4092 -744 4138 -732
rect 4188 -740 4234 -732
rect 4092 -972 4098 -744
rect 4132 -972 4138 -744
rect 4092 -984 4138 -972
rect 4182 -744 4240 -740
rect 4182 -752 4194 -744
rect 4228 -752 4240 -744
rect 4238 -980 4240 -752
rect 4098 -1110 4132 -984
rect 4182 -992 4240 -980
rect 4284 -744 4330 -732
rect 4380 -740 4426 -732
rect 4284 -972 4290 -744
rect 4324 -972 4330 -744
rect 4284 -984 4330 -972
rect 4374 -744 4432 -740
rect 4374 -752 4386 -744
rect 4420 -752 4432 -744
rect 4374 -980 4376 -752
rect 4290 -1110 4324 -984
rect 4374 -992 4432 -980
rect 4476 -744 4522 -732
rect 4572 -740 4618 -732
rect 4476 -972 4482 -744
rect 4516 -972 4522 -744
rect 4476 -984 4522 -972
rect 4566 -744 4624 -740
rect 4566 -752 4578 -744
rect 4612 -752 4624 -744
rect 4566 -980 4568 -752
rect 4482 -1110 4516 -984
rect 4566 -992 4624 -980
rect 4668 -744 4714 -732
rect 4764 -740 4810 -732
rect 4668 -972 4674 -744
rect 4708 -972 4714 -744
rect 4668 -984 4714 -972
rect 4758 -744 4816 -740
rect 4758 -752 4770 -744
rect 4804 -752 4816 -744
rect 4814 -980 4816 -752
rect 4674 -1110 4708 -984
rect 4758 -992 4816 -980
rect 4860 -744 4906 -732
rect 4956 -742 5002 -732
rect 4860 -972 4866 -744
rect 4900 -972 4906 -744
rect 4860 -984 4906 -972
rect 4950 -744 5008 -742
rect 4950 -752 4962 -744
rect 4996 -752 5008 -744
rect 5006 -980 5008 -752
rect 4866 -1110 4900 -984
rect 4950 -994 5008 -980
rect 5052 -744 5098 -732
rect 5148 -742 5194 -732
rect 5052 -972 5058 -744
rect 5092 -972 5098 -744
rect 5052 -984 5098 -972
rect 5144 -744 5202 -742
rect 5144 -752 5154 -744
rect 5188 -752 5202 -744
rect 5200 -980 5202 -752
rect 5058 -1110 5092 -984
rect 5144 -994 5202 -980
rect 5244 -744 5290 -732
rect 5340 -740 5386 -732
rect 5244 -972 5250 -744
rect 5284 -972 5290 -744
rect 5244 -984 5290 -972
rect 5334 -744 5392 -740
rect 5334 -752 5346 -744
rect 5380 -752 5392 -744
rect 5334 -980 5336 -752
rect 5250 -1110 5284 -984
rect 5334 -992 5392 -980
rect 5436 -744 5482 -732
rect 5532 -740 5578 -732
rect 5436 -972 5442 -744
rect 5476 -972 5482 -744
rect 5436 -984 5482 -972
rect 5526 -744 5584 -740
rect 5526 -752 5538 -744
rect 5572 -752 5584 -744
rect 5582 -980 5584 -752
rect 5442 -1110 5476 -984
rect 5526 -992 5584 -980
rect 5628 -744 5674 -732
rect 5724 -740 5770 -732
rect 5628 -972 5634 -744
rect 5668 -972 5674 -744
rect 5628 -984 5674 -972
rect 5718 -744 5776 -740
rect 5718 -752 5730 -744
rect 5764 -752 5776 -744
rect 5774 -980 5776 -752
rect 5634 -1110 5668 -984
rect 5718 -992 5776 -980
rect 5820 -744 5866 -732
rect 5916 -742 5964 -732
rect 5820 -972 5826 -744
rect 5860 -972 5866 -744
rect 5820 -984 5866 -972
rect 5910 -744 5970 -742
rect 5910 -752 5922 -744
rect 5956 -752 5970 -744
rect 5910 -980 5912 -752
rect 5968 -980 5970 -752
rect 5835 -1110 5865 -984
rect 5910 -992 5970 -980
rect -278 -1140 5865 -1110
rect -278 -1142 5864 -1140
rect -404 -1218 1666 -1216
rect -404 -1314 5988 -1218
rect -404 -1320 1462 -1314
rect -404 -1398 -326 -1320
rect -398 -1708 -326 -1398
rect 5970 -1708 5988 -1314
rect -398 -1832 5988 -1708
<< via1 >>
rect -188 766 5906 1208
rect 502 506 558 508
rect 502 278 510 506
rect 510 278 544 506
rect 544 278 558 506
rect 502 276 558 278
rect 696 278 710 506
rect 710 278 746 506
rect 746 278 756 506
rect -170 180 28 186
rect -170 136 28 180
rect -170 132 28 136
rect 0 10 54 70
rect 900 282 956 506
rect 1100 280 1156 508
rect 1302 280 1358 508
rect 1502 280 1558 508
rect 1934 326 1990 556
rect 2126 326 2180 554
rect 2340 326 2396 554
rect 200 12 254 72
rect 500 10 510 70
rect 510 10 544 70
rect 544 10 554 70
rect 700 10 710 70
rect 710 10 744 70
rect 744 10 754 70
rect 900 10 952 70
rect 1100 12 1152 72
rect 1304 10 1356 70
rect 1504 12 1556 72
rect 354 -86 772 -78
rect 354 -122 770 -86
rect 770 -122 772 -86
rect 354 -130 772 -122
rect 1930 14 1986 74
rect 2534 326 2590 554
rect 2724 326 2780 554
rect 2918 324 2974 552
rect 3110 326 3166 554
rect 2122 14 2178 74
rect 2344 14 2398 74
rect 2536 14 2590 74
rect 2728 14 2782 74
rect 2920 14 2974 74
rect 3114 14 3168 74
rect 40 -412 96 -408
rect 40 -460 48 -412
rect 48 -460 86 -412
rect 86 -460 96 -412
rect 202 -406 254 -404
rect 202 -466 210 -406
rect 210 -466 244 -406
rect 244 -466 254 -406
rect 202 -468 254 -466
rect 502 -464 510 -404
rect 510 -464 544 -404
rect 544 -464 554 -404
rect 702 -464 710 -404
rect 710 -464 744 -404
rect 744 -464 754 -404
rect 906 -468 916 -408
rect 916 -468 950 -408
rect 950 -468 958 -408
rect -40 -534 274 -526
rect -40 -576 272 -534
rect 272 -576 274 -534
rect -40 -584 274 -576
rect 1106 -470 1116 -410
rect 1116 -470 1150 -410
rect 1150 -470 1158 -410
rect 1310 -468 1318 -408
rect 1318 -468 1352 -408
rect 1352 -468 1362 -408
rect 1510 -470 1518 -410
rect 1518 -470 1552 -410
rect 1552 -470 1562 -410
rect 1930 -470 1940 -410
rect 1940 -470 1974 -410
rect 1974 -470 1986 -410
rect 2122 -470 2132 -410
rect 2132 -470 2166 -410
rect 2166 -470 2178 -410
rect 2344 -470 2354 -410
rect 2354 -470 2388 -410
rect 2388 -470 2398 -410
rect 2536 -470 2546 -410
rect 2546 -470 2580 -410
rect 2580 -470 2590 -410
rect 2728 -470 2738 -410
rect 2738 -470 2772 -410
rect 2772 -470 2782 -410
rect 2920 -470 2930 -410
rect 2930 -470 2964 -410
rect 2964 -470 2974 -410
rect 3114 -470 3122 -410
rect 3122 -470 3156 -410
rect 3156 -470 3168 -410
rect 502 -900 510 -696
rect 510 -900 544 -696
rect 544 -900 554 -696
rect 700 -900 710 -696
rect 710 -900 744 -696
rect 744 -900 752 -696
rect 906 -904 916 -680
rect 916 -904 950 -680
rect 950 -904 962 -680
rect 1106 -906 1116 -678
rect 1116 -906 1150 -678
rect 1150 -906 1162 -678
rect 1308 -906 1318 -678
rect 1318 -906 1352 -678
rect 1352 -906 1364 -678
rect 1698 -576 1858 -522
rect 3416 -470 3426 -410
rect 3426 -470 3460 -410
rect 3460 -470 3472 -410
rect 3608 -470 3618 -410
rect 3618 -470 3652 -410
rect 3652 -470 3664 -410
rect 3798 -470 3810 -410
rect 3810 -470 3844 -410
rect 3844 -470 3854 -410
rect 3990 -470 4002 -410
rect 4002 -470 4036 -410
rect 4036 -470 4046 -410
rect 4182 -470 4194 -410
rect 4194 -470 4228 -410
rect 4228 -470 4238 -410
rect 4374 -470 4386 -410
rect 4386 -470 4420 -410
rect 4420 -470 4430 -410
rect 4566 -470 4578 -410
rect 4578 -470 4612 -410
rect 4612 -470 4622 -410
rect 4760 -470 4770 -410
rect 4770 -470 4804 -410
rect 4804 -470 4816 -410
rect 4952 -470 4962 -410
rect 4962 -470 4996 -410
rect 4996 -470 5008 -410
rect 5142 -470 5154 -410
rect 5154 -470 5188 -410
rect 5188 -470 5198 -410
rect 5336 -470 5346 -410
rect 5346 -470 5380 -410
rect 5380 -470 5392 -410
rect 5526 -470 5538 -410
rect 5538 -470 5572 -410
rect 5572 -470 5582 -410
rect 5718 -470 5730 -410
rect 5730 -470 5764 -410
rect 5764 -470 5774 -410
rect 5910 -470 5922 -410
rect 5922 -470 5956 -410
rect 5956 -470 5966 -410
rect 1508 -906 1518 -678
rect 1518 -906 1552 -678
rect 1552 -906 1564 -678
rect 1934 -950 1944 -722
rect 1944 -950 1978 -722
rect 1978 -950 1990 -722
rect 1934 -952 1990 -950
rect 2126 -950 2136 -722
rect 2136 -950 2170 -722
rect 2170 -950 2180 -722
rect 2340 -950 2352 -722
rect 2352 -950 2386 -722
rect 2386 -950 2396 -722
rect 2534 -950 2544 -722
rect 2544 -950 2578 -722
rect 2578 -950 2590 -722
rect 2724 -950 2736 -722
rect 2736 -950 2770 -722
rect 2770 -950 2780 -722
rect 2918 -722 2974 -720
rect 2918 -948 2928 -722
rect 2928 -948 2962 -722
rect 2962 -948 2974 -722
rect 3110 -950 3120 -722
rect 3120 -950 3154 -722
rect 3154 -950 3166 -722
rect 3414 -972 3426 -752
rect 3426 -972 3460 -752
rect 3460 -972 3470 -752
rect 3414 -980 3470 -972
rect 3606 -972 3618 -752
rect 3618 -972 3652 -752
rect 3652 -972 3662 -752
rect 3606 -980 3662 -972
rect 3800 -972 3810 -752
rect 3810 -972 3844 -752
rect 3844 -972 3856 -752
rect 3800 -980 3856 -972
rect 3992 -972 4002 -752
rect 4002 -972 4036 -752
rect 4036 -972 4048 -752
rect 3992 -980 4048 -972
rect 4182 -972 4194 -752
rect 4194 -972 4228 -752
rect 4228 -972 4238 -752
rect 4182 -980 4238 -972
rect 4376 -972 4386 -752
rect 4386 -972 4420 -752
rect 4420 -972 4432 -752
rect 4376 -980 4432 -972
rect 4568 -972 4578 -752
rect 4578 -972 4612 -752
rect 4612 -972 4624 -752
rect 4568 -980 4624 -972
rect 4758 -972 4770 -752
rect 4770 -972 4804 -752
rect 4804 -972 4814 -752
rect 4758 -980 4814 -972
rect 4950 -972 4962 -752
rect 4962 -972 4996 -752
rect 4996 -972 5006 -752
rect 4950 -980 5006 -972
rect 5144 -972 5154 -752
rect 5154 -972 5188 -752
rect 5188 -972 5200 -752
rect 5144 -980 5200 -972
rect 5336 -972 5346 -752
rect 5346 -972 5380 -752
rect 5380 -972 5392 -752
rect 5336 -980 5392 -972
rect 5526 -972 5538 -752
rect 5538 -972 5572 -752
rect 5572 -972 5582 -752
rect 5526 -980 5582 -972
rect 5718 -972 5730 -752
rect 5730 -972 5764 -752
rect 5764 -972 5774 -752
rect 5718 -980 5774 -972
rect 5912 -972 5922 -752
rect 5922 -972 5956 -752
rect 5956 -972 5968 -752
rect 5912 -980 5968 -972
rect 1462 -1320 5970 -1314
rect -326 -1708 5970 -1320
<< metal2 >>
rect -280 1208 6008 1268
rect -280 766 -188 1208
rect 5906 766 6008 1208
rect -280 698 6008 766
rect 1924 556 2002 568
rect 488 508 566 518
rect 488 276 502 508
rect 558 276 566 508
rect 488 266 566 276
rect 680 506 768 518
rect 680 278 696 506
rect 756 278 768 506
rect 680 264 768 278
rect 890 506 966 522
rect 890 282 900 506
rect 956 282 966 506
rect 890 266 966 282
rect 1088 508 1160 524
rect 1088 280 1100 508
rect 1156 280 1160 508
rect 1088 268 1160 280
rect 1290 508 1362 522
rect 1290 280 1302 508
rect 1358 280 1362 508
rect 1290 266 1362 280
rect 1490 508 1562 522
rect 1490 280 1502 508
rect 1558 280 1562 508
rect 1924 326 1934 556
rect 1990 326 2002 556
rect 1924 314 2002 326
rect 2114 556 2192 566
rect 2114 326 2126 556
rect 2182 326 2192 556
rect 2114 312 2192 326
rect 2332 554 2404 566
rect 2332 326 2340 554
rect 2396 326 2404 554
rect 2332 312 2404 326
rect 2528 554 2600 564
rect 2528 326 2534 554
rect 2590 326 2600 554
rect 2528 314 2600 326
rect 2718 554 2790 566
rect 2718 326 2724 554
rect 2780 326 2790 554
rect 2718 316 2790 326
rect 2912 552 2984 564
rect 2912 324 2918 552
rect 2974 324 2984 552
rect 2912 314 2984 324
rect 3100 554 3172 566
rect 3100 326 3110 554
rect 3166 326 3172 554
rect 3100 316 3172 326
rect 1490 266 1562 280
rect -182 190 40 198
rect -182 128 -170 190
rect 28 128 40 190
rect -182 120 40 128
rect 3136 86 3452 88
rect 1506 84 3452 86
rect -2 80 56 82
rect 202 80 252 82
rect 818 80 3452 84
rect -2 74 3452 80
rect -2 72 1930 74
rect -2 70 200 72
rect -2 10 0 70
rect 54 12 200 70
rect 254 70 1100 72
rect 254 12 500 70
rect 54 10 500 12
rect 554 10 700 70
rect 754 10 900 70
rect 952 12 1100 70
rect 1152 70 1504 72
rect 1152 12 1304 70
rect 952 10 1304 12
rect 1356 12 1504 70
rect 1556 14 1930 72
rect 1986 14 2122 74
rect 2178 14 2344 74
rect 2398 14 2536 74
rect 2590 14 2728 74
rect 2782 14 2920 74
rect 2974 14 3114 74
rect 3168 14 3452 74
rect 1556 12 3452 14
rect 1356 10 3452 12
rect -2 -2 3452 10
rect 202 -262 252 -2
rect 1506 -4 3452 -2
rect 3136 -6 3452 -4
rect 338 -74 792 -66
rect 338 -132 354 -74
rect 774 -132 792 -74
rect -398 -264 -284 -262
rect 146 -264 254 -262
rect -398 -322 254 -264
rect -398 -1216 -322 -322
rect 32 -388 100 -322
rect 32 -408 102 -388
rect 202 -398 252 -322
rect 1476 -396 3184 -392
rect 840 -398 3184 -396
rect 32 -460 40 -408
rect 96 -460 102 -408
rect 32 -486 102 -460
rect 190 -404 5968 -398
rect 190 -468 202 -404
rect 254 -464 502 -404
rect 554 -464 702 -404
rect 754 -408 5968 -404
rect 754 -464 906 -408
rect 254 -468 906 -464
rect 958 -410 1310 -408
rect 958 -468 1106 -410
rect 190 -470 1106 -468
rect 1158 -468 1310 -410
rect 1362 -410 5968 -408
rect 1362 -468 1510 -410
rect 1158 -470 1510 -468
rect 1562 -470 1930 -410
rect 1986 -470 2122 -410
rect 2178 -470 2344 -410
rect 2398 -470 2536 -410
rect 2590 -470 2728 -410
rect 2782 -470 2920 -410
rect 2974 -470 3114 -410
rect 3168 -470 3416 -410
rect 3472 -470 3608 -410
rect 3664 -470 3798 -410
rect 3854 -470 3990 -410
rect 4046 -470 4182 -410
rect 4238 -470 4374 -410
rect 4430 -470 4566 -410
rect 4622 -470 4760 -410
rect 4816 -470 4952 -410
rect 5008 -470 5142 -410
rect 5198 -470 5336 -410
rect 5392 -470 5526 -410
rect 5582 -470 5718 -410
rect 5774 -470 5910 -410
rect 5966 -470 5968 -410
rect 190 -478 5968 -470
rect 202 -480 252 -478
rect 840 -482 5968 -478
rect 840 -484 912 -482
rect 1476 -484 1980 -482
rect 3380 -484 5968 -482
rect -56 -526 286 -516
rect -56 -584 -40 -526
rect 274 -584 286 -526
rect 1682 -520 1872 -518
rect 1682 -576 1698 -520
rect 1858 -576 1872 -520
rect 1682 -578 1872 -576
rect -56 -592 286 -584
rect 896 -680 972 -664
rect 494 -696 566 -684
rect 494 -900 502 -696
rect 558 -900 566 -696
rect 494 -912 566 -900
rect 696 -696 768 -684
rect 696 -900 700 -696
rect 756 -900 768 -696
rect 696 -912 768 -900
rect 896 -904 906 -680
rect 962 -904 972 -680
rect 896 -920 972 -904
rect 1094 -678 1166 -666
rect 1094 -906 1106 -678
rect 1162 -906 1166 -678
rect 1094 -922 1166 -906
rect 1296 -678 1368 -664
rect 1296 -906 1308 -678
rect 1364 -906 1368 -678
rect 1296 -920 1368 -906
rect 1496 -678 1568 -664
rect 1496 -906 1508 -678
rect 1564 -906 1568 -678
rect 1496 -920 1568 -906
rect 1924 -722 2002 -710
rect 1924 -952 1934 -722
rect 1990 -952 2002 -722
rect 1924 -964 2002 -952
rect 2114 -722 2192 -708
rect 2114 -952 2126 -722
rect 2182 -952 2192 -722
rect 2114 -962 2192 -952
rect 2332 -722 2404 -708
rect 2332 -950 2340 -722
rect 2396 -950 2404 -722
rect 2332 -962 2404 -950
rect 2528 -722 2600 -710
rect 2528 -950 2534 -722
rect 2590 -950 2600 -722
rect 2528 -960 2600 -950
rect 2718 -722 2790 -712
rect 2718 -950 2724 -722
rect 2780 -950 2790 -722
rect 2718 -962 2790 -950
rect 2912 -720 2984 -710
rect 2912 -948 2918 -720
rect 2974 -948 2984 -720
rect 2912 -960 2984 -948
rect 3100 -722 3172 -712
rect 3100 -950 3110 -722
rect 3166 -950 3172 -722
rect 3100 -962 3172 -950
rect 3374 -752 5968 -740
rect 3374 -980 3414 -752
rect 3470 -980 3606 -752
rect 3662 -980 3800 -752
rect 3856 -980 3992 -752
rect 4048 -980 4182 -752
rect 4238 -980 4376 -752
rect 4432 -980 4568 -752
rect 4624 -980 4758 -752
rect 4814 -980 4950 -752
rect 5006 -980 5144 -752
rect 5200 -980 5336 -752
rect 5392 -980 5526 -752
rect 5582 -980 5718 -752
rect 5774 -980 5912 -752
rect 3374 -992 5968 -980
rect -404 -1218 1666 -1216
rect -404 -1314 5988 -1218
rect -404 -1320 1462 -1314
rect -404 -1398 -326 -1320
rect -400 -1708 -326 -1398
rect 5970 -1708 5988 -1314
rect -400 -1716 -320 -1708
rect 1250 -1716 5988 -1708
rect -400 -1826 5988 -1716
rect -398 -1832 5988 -1826
<< via2 >>
rect -188 766 5906 1208
rect 502 276 558 508
rect 696 278 756 506
rect 900 282 956 506
rect 1100 280 1156 508
rect 1302 280 1358 508
rect 1502 280 1558 508
rect 1934 326 1990 556
rect 2126 554 2182 556
rect 2126 326 2180 554
rect 2180 326 2182 554
rect 2340 326 2396 554
rect 2534 326 2590 554
rect 2724 326 2780 554
rect 2918 324 2974 552
rect 3110 326 3166 554
rect -170 186 28 190
rect -170 132 28 186
rect -170 128 28 132
rect 354 -78 774 -74
rect 354 -130 772 -78
rect 772 -130 774 -78
rect 354 -132 774 -130
rect -40 -584 274 -526
rect 1698 -522 1858 -520
rect 1698 -576 1858 -522
rect 502 -900 554 -696
rect 554 -900 558 -696
rect 700 -900 752 -696
rect 752 -900 756 -696
rect 906 -904 962 -680
rect 1106 -906 1162 -678
rect 1308 -906 1364 -678
rect 1508 -906 1564 -678
rect 1934 -952 1990 -722
rect 2126 -950 2180 -722
rect 2180 -950 2182 -722
rect 2126 -952 2182 -950
rect 2340 -950 2396 -722
rect 2534 -950 2590 -722
rect 2724 -950 2780 -722
rect 2918 -948 2974 -720
rect 3110 -950 3166 -722
rect 1462 -1320 5970 -1314
rect -326 -1708 5970 -1320
rect -320 -1716 1250 -1708
<< metal3 >>
rect -284 1208 6010 1274
rect -284 766 -188 1208
rect 5906 766 6010 1208
rect -284 698 6010 766
rect 1924 566 2002 568
rect 2120 566 3190 570
rect 1924 556 3190 566
rect 486 508 1576 518
rect 486 276 502 508
rect 558 506 1100 508
rect 558 278 696 506
rect 756 282 900 506
rect 956 282 1100 506
rect 756 280 1100 282
rect 1156 280 1302 508
rect 1358 280 1502 508
rect 1558 280 1576 508
rect 1924 326 1934 556
rect 1990 326 2126 556
rect 2182 554 3190 556
rect 2182 326 2340 554
rect 2396 326 2534 554
rect 2590 326 2724 554
rect 2780 552 3110 554
rect 2780 326 2918 552
rect 1924 324 2918 326
rect 2974 326 3110 552
rect 3166 326 3190 554
rect 2974 324 3190 326
rect 1924 314 3190 324
rect 2114 312 3190 314
rect 756 278 1576 280
rect 558 276 1576 278
rect 486 266 1576 276
rect 680 264 768 266
rect -196 190 40 198
rect -196 128 -170 190
rect 28 128 40 190
rect -196 120 40 128
rect -196 -522 -124 120
rect 338 -69 792 -66
rect 338 -74 1817 -69
rect 338 -132 354 -74
rect 774 -132 1817 -74
rect 338 -135 1817 -132
rect 338 -140 792 -135
rect 1751 -510 1817 -135
rect -56 -522 286 -516
rect -196 -526 286 -522
rect -196 -584 -40 -526
rect 274 -584 286 -526
rect -196 -592 286 -584
rect 1682 -520 1874 -510
rect 1682 -576 1698 -520
rect 1858 -576 1874 -520
rect 1682 -586 1874 -576
rect -196 -594 224 -592
rect 1751 -599 1817 -586
rect 654 -678 1582 -664
rect 654 -680 1106 -678
rect 654 -686 906 -680
rect 486 -696 906 -686
rect 486 -900 502 -696
rect 558 -900 700 -696
rect 756 -900 906 -696
rect 486 -904 906 -900
rect 962 -904 1106 -680
rect 486 -906 1106 -904
rect 1162 -906 1308 -678
rect 1364 -906 1508 -678
rect 1564 -906 1582 -678
rect 486 -914 1582 -906
rect 654 -916 1582 -914
rect 1922 -720 3190 -708
rect 1922 -722 2918 -720
rect 1922 -952 1934 -722
rect 1990 -952 2126 -722
rect 2182 -950 2340 -722
rect 2396 -950 2534 -722
rect 2590 -950 2724 -722
rect 2780 -948 2918 -722
rect 2974 -722 3190 -720
rect 2974 -948 3110 -722
rect 2780 -950 3110 -948
rect 3166 -950 3190 -722
rect 2182 -952 3190 -950
rect 1922 -966 3190 -952
rect -404 -1218 1666 -1216
rect -404 -1314 5988 -1218
rect -404 -1320 1462 -1314
rect -404 -1398 -326 -1320
rect -400 -1708 -326 -1398
rect 5970 -1708 5988 -1314
rect -400 -1716 -320 -1708
rect 1250 -1716 5988 -1708
rect -400 -1826 5988 -1716
rect -398 -1832 5988 -1826
<< via3 >>
rect -188 766 5906 1208
rect 1462 -1320 5970 -1314
rect -326 -1708 5970 -1320
rect -320 -1716 1250 -1708
<< metal4 >>
rect 1328 1254 6012 1266
rect -284 1208 6012 1254
rect -284 840 -188 1208
rect -280 766 -188 840
rect 5906 766 6012 1208
rect -280 678 6012 766
rect 864 676 1416 678
rect -404 -1218 1666 -1216
rect -404 -1314 5988 -1218
rect -404 -1320 1462 -1314
rect -404 -1398 -326 -1320
rect -400 -1708 -326 -1398
rect 5970 -1708 5988 -1314
rect -400 -1716 -320 -1708
rect 1250 -1716 5988 -1708
rect -400 -1826 5988 -1716
rect -398 -1832 5988 -1826
<< via4 >>
rect 1462 -1320 5970 -1314
rect -326 -1708 5970 -1320
rect -320 -1716 1250 -1708
<< metal5 >>
rect -404 -1314 5994 -1216
rect -404 -1320 1462 -1314
rect -404 -1322 -326 -1320
rect -410 -1708 -326 -1322
rect 5970 -1708 5994 -1314
rect -410 -1716 -320 -1708
rect 1250 -1716 5994 -1708
rect -410 -1830 5994 -1716
rect -410 -1832 5988 -1830
use inverter_27x  inverter_27x_0 ~/Desktop/charge_pumps2/layout_files
timestamp 1698771642
transform 1 0 4518 0 1 -1396
box -1236 1310 1512 2140
use sky130_fd_pr__nfet_01v8_5ACVEW  sky130_fd_pr__nfet_01v8_5ACVEW_0 ~/Desktop/charge_pumps2/layout_files
timestamp 1698771642
transform 1 0 2101 0 1 44
box -173 -130 173 130
use sky130_fd_pr__nfet_01v8_D4CDWR  sky130_fd_pr__nfet_01v8_D4CDWR_0 ~/Desktop/charge_pumps2/layout_files
timestamp 1698771642
transform 1 0 2803 0 1 44
box -461 -130 461 130
use sky130_fd_pr__nfet_01v8_DQBD8A  sky130_fd_pr__nfet_01v8_DQBD8A_0 ~/Desktop/charge_pumps2/layout_files
timestamp 1698771642
transform 1 0 971 0 1 40
box -73 -68 73 68
use sky130_fd_pr__nfet_01v8_DQBD8A  sky130_fd_pr__nfet_01v8_DQBD8A_1
timestamp 1698771642
transform 1 0 1171 0 1 42
box -73 -68 73 68
use sky130_fd_pr__nfet_01v8_DQBD8A  sky130_fd_pr__nfet_01v8_DQBD8A_2
timestamp 1698771642
transform 1 0 1373 0 1 40
box -73 -68 73 68
use sky130_fd_pr__nfet_01v8_DQBD8A  sky130_fd_pr__nfet_01v8_DQBD8A_3
timestamp 1698771642
transform 1 0 1573 0 1 42
box -73 -68 73 68
use sky130_fd_pr__nfet_01v8_KMMFCM  sky130_fd_pr__nfet_01v8_KMMFCM_0 ~/Desktop/charge_pumps2/layout_files
timestamp 1698771642
transform 1 0 71 0 1 40
box -73 -68 73 68
use sky130_fd_pr__nfet_01v8_KMMFCM  sky130_fd_pr__nfet_01v8_KMMFCM_1
timestamp 1698771642
transform 1 0 359 0 1 42
box -73 -68 73 68
use sky130_fd_pr__nfet_01v8_KMMFCM  sky130_fd_pr__nfet_01v8_KMMFCM_2
timestamp 1698771642
transform 1 0 271 0 1 42
box -73 -68 73 68
use sky130_fd_pr__pfet_01v8_29EZRJ  sky130_fd_pr__pfet_01v8_29EZRJ_0 ~/Desktop/charge_pumps2/layout_files
timestamp 1698771642
transform 1 0 71 0 1 392
box -109 -188 109 188
use sky130_fd_pr__pfet_01v8_29EZRJ  sky130_fd_pr__pfet_01v8_29EZRJ_1
timestamp 1698771642
transform 1 0 359 0 1 440
box -109 -188 109 188
use sky130_fd_pr__pfet_01v8_29EZRJ  sky130_fd_pr__pfet_01v8_29EZRJ_2
timestamp 1698771642
transform 1 0 271 0 1 440
box -109 -188 109 188
use sky130_fd_pr__pfet_01v8_29EZRJ  sky130_fd_pr__pfet_01v8_29EZRJ_3
timestamp 1698771642
transform 1 0 971 0 1 394
box -109 -188 109 188
use sky130_fd_pr__pfet_01v8_FBZ64Q  sky130_fd_pr__pfet_01v8_FBZ64Q_0 ~/Desktop/charge_pumps2/layout_files
timestamp 1698771642
transform 1 0 2801 0 1 440
box -497 -226 497 226
use sky130_fd_pr__pfet_01v8_FL984Q  sky130_fd_pr__pfet_01v8_FL984Q_0 ~/Desktop/charge_pumps2/layout_files
timestamp 1698771642
transform 1 0 2105 0 1 440
box -209 -226 209 226
use sky130_fd_pr__pfet_01v8_FXZ64Q  sky130_fd_pr__pfet_01v8_FXZ64Q_0 ~/Desktop/charge_pumps2/layout_files
timestamp 1698771642
transform 1 0 1171 0 1 394
box -109 -188 109 188
use sky130_fd_pr__pfet_01v8_FXZ64Q  sky130_fd_pr__pfet_01v8_FXZ64Q_1
timestamp 1698771642
transform 1 0 1373 0 1 394
box -109 -188 109 188
use sky130_fd_pr__pfet_01v8_FXZ64Q  sky130_fd_pr__pfet_01v8_FXZ64Q_2
timestamp 1698771642
transform 1 0 1573 0 1 394
box -109 -188 109 188
<< labels >>
rlabel metal3 -172 -142 -172 -142 1 clk_in
port 1 n
rlabel via3 4264 1018 4264 1018 1 vdd
port 2 n
rlabel via4 5274 -1522 5274 -1522 1 gnd
port 3 n
rlabel metal1 5976 -124 5976 -124 1 clk
port 4 n
rlabel metal1 5794 -262 5794 -262 1 clkb
port 5 n
<< end >>
