magic
tech sky130A
magscale 1 2
timestamp 1698914177
<< psubdiff >>
rect 5661 -409 5748 -383
rect 5661 -450 5688 -409
rect 5722 -450 5748 -409
rect 5661 -475 5748 -450
<< psubdiffcont >>
rect 5688 -450 5722 -409
<< poly >>
rect 38 -356 173 -322
rect 38 -375 72 -356
rect 932 -359 1061 -329
rect 932 -402 962 -359
rect 1890 -362 2013 -332
rect 2848 -352 2977 -322
rect 3830 -329 3860 -324
rect 1890 -394 1920 -362
rect 2848 -384 2878 -352
rect 3830 -359 3959 -329
rect 4772 -356 4901 -326
rect 3830 -386 3860 -359
rect 4772 -388 4802 -356
<< locali >>
rect 302 -290 988 -258
rect 5661 -409 5748 -383
rect 5661 -451 5687 -409
rect 5722 -451 5748 -409
rect 5661 -475 5748 -451
rect -16 -612 5796 -526
rect -16 -614 666 -612
<< viali >>
rect 5687 -450 5688 -409
rect 5688 -450 5722 -409
rect 5687 -451 5722 -450
<< metal1 >>
rect -224 1534 6008 1598
rect -242 1330 -232 1534
rect 5994 1465 6008 1534
rect 5994 1423 6876 1465
rect 5994 1330 6008 1423
rect -224 1244 6008 1330
rect 424 1064 528 1244
rect 5503 1228 5623 1244
rect 5740 1217 5856 1244
rect -274 960 914 1064
rect -660 465 -344 466
rect -1681 458 -344 465
rect -1681 399 -636 458
rect -1476 -858 -1408 -842
rect -1476 -984 -1466 -858
rect -1412 -984 -1408 -858
rect -1240 -878 -1190 -846
rect -1476 -1000 -1408 -984
rect -855 -1171 -789 399
rect -660 398 -636 399
rect -374 398 -344 458
rect -660 384 -344 398
rect -274 -578 -170 960
rect 424 930 528 960
rect 2438 884 2524 896
rect 2436 828 2446 884
rect 2508 828 2524 884
rect 2438 824 2524 828
rect 870 244 974 258
rect 870 190 882 244
rect 954 190 974 244
rect 1254 192 1264 250
rect 1346 192 1356 250
rect 2424 192 2434 252
rect 2508 192 2518 252
rect 2812 190 2822 248
rect 2892 190 2902 248
rect 870 188 974 190
rect 6068 -88 6448 -78
rect 6068 -144 6090 -88
rect 6428 -144 6448 -88
rect 6068 -154 6448 -144
rect -12 -432 16 -212
rect 302 -290 988 -264
rect 124 -360 740 -326
rect 882 -420 916 -290
rect 1014 -376 1646 -326
rect 1840 -416 1874 -260
rect 1968 -372 2600 -322
rect -14 -460 790 -432
rect -12 -470 16 -460
rect 878 -472 1680 -420
rect 1840 -454 2646 -416
rect 1844 -468 2646 -454
rect 2794 -424 2828 -260
rect 2934 -372 3560 -330
rect 3780 -424 3814 -266
rect 3920 -376 4546 -334
rect 4722 -420 4756 -274
rect 4854 -374 5480 -332
rect 5680 -397 5728 -213
rect 5680 -409 5730 -397
rect 2794 -476 3596 -424
rect 3778 -476 4580 -424
rect 4720 -472 5522 -420
rect 5680 -451 5687 -409
rect 5722 -451 5730 -409
rect 5680 -464 5730 -451
rect 26 -520 664 -516
rect -16 -526 666 -520
rect -16 -578 5796 -526
rect -274 -612 5796 -578
rect -274 -614 666 -612
rect -274 -682 2 -614
rect -506 -1162 -416 -1160
rect -506 -1171 -190 -1162
rect -855 -1176 -190 -1171
rect -855 -1232 -440 -1176
rect -224 -1232 -190 -1176
rect -855 -1237 -190 -1232
rect -506 -1244 -190 -1237
rect -478 -1246 -190 -1244
rect -618 -1444 -244 -1420
rect 826 -1442 836 -1378
rect 926 -1442 936 -1378
rect 1212 -1440 1222 -1376
rect 1312 -1440 1322 -1376
rect 2366 -1386 2480 -1372
rect 2366 -1442 2404 -1386
rect 2472 -1442 2482 -1386
rect 2366 -1444 2480 -1442
rect 2778 -1444 2788 -1390
rect 2852 -1444 2862 -1390
rect -754 -1518 -716 -1514
rect -754 -1546 -656 -1518
rect -618 -1522 -572 -1444
rect -294 -1522 -244 -1444
rect -754 -1590 -716 -1546
rect -618 -1548 -244 -1522
rect -170 -1820 5588 -1818
rect 5864 -1820 5962 -178
rect 6073 -846 6111 -154
rect 6834 -580 6876 1423
rect 8464 -806 8653 -756
rect 6073 -884 6239 -846
rect 6074 -966 6242 -930
rect 6074 -1700 6110 -966
rect 6834 -1084 6876 -1082
rect 6830 -1124 6876 -1084
rect 6070 -1708 6440 -1700
rect 6070 -1712 6094 -1708
rect 6408 -1712 6440 -1708
rect 6070 -1770 6092 -1712
rect 6434 -1770 6440 -1712
rect 6070 -1780 6440 -1770
rect -170 -1890 6052 -1820
rect -146 -1936 6052 -1890
rect -154 -2114 -144 -1936
rect 6022 -2048 6052 -1936
rect 6830 -2048 6866 -1124
rect 6022 -2084 6866 -2048
rect 6022 -2114 6052 -2084
rect -146 -2214 6052 -2114
<< via1 >>
rect -232 1330 5994 1534
rect -1466 -984 -1412 -858
rect -636 398 -374 458
rect 2446 828 2508 884
rect 882 190 954 244
rect 1264 192 1346 250
rect 2434 192 2508 252
rect 2822 190 2892 248
rect 6090 -144 6428 -88
rect -440 -1232 -224 -1176
rect 836 -1442 926 -1378
rect 1222 -1440 1312 -1376
rect 2404 -1442 2472 -1386
rect 2788 -1444 2852 -1390
rect -572 -1522 -294 -1444
rect 6094 -1712 6408 -1708
rect 6092 -1770 6434 -1712
rect -144 -2114 6022 -1936
<< metal2 >>
rect -232 1534 5994 1544
rect -232 1320 5994 1330
rect 2438 884 2524 896
rect 2438 828 2446 884
rect 2508 828 2524 884
rect 2438 824 2524 828
rect 2446 818 2508 824
rect -660 458 -344 466
rect -660 398 -636 458
rect -374 398 -344 458
rect -660 384 -344 398
rect -1681 296 1314 326
rect -1476 -858 -1408 -842
rect -1476 -984 -1470 -858
rect -1412 -984 -1408 -858
rect -1476 -1000 -1408 -984
rect -701 -1286 -671 296
rect 1284 262 1314 296
rect -642 238 -302 246
rect -642 160 -608 238
rect -328 224 -302 238
rect 870 244 974 258
rect 870 224 882 244
rect -328 190 882 224
rect 954 190 974 244
rect 1258 250 1358 262
rect 1258 192 1264 250
rect 1346 192 1358 250
rect 1258 190 1358 192
rect 2434 252 2508 262
rect -328 188 974 190
rect -328 160 -302 188
rect 882 180 954 188
rect 1264 182 1346 190
rect 2434 182 2508 192
rect 2822 248 2892 258
rect 2822 180 2892 190
rect -642 140 -302 160
rect 4746 -80 4874 -70
rect 6068 -88 6448 -78
rect 6068 -144 6090 -88
rect 6428 -144 6448 -88
rect 6068 -154 6448 -144
rect 4746 -166 4874 -156
rect 2764 -732 2872 -722
rect 2764 -808 2872 -798
rect -478 -1176 -190 -1162
rect -478 -1232 -440 -1176
rect -224 -1232 -190 -1176
rect -478 -1246 -190 -1232
rect -701 -1318 1284 -1286
rect -701 -1351 -671 -1318
rect 776 -1366 954 -1364
rect 1252 -1366 1284 -1318
rect 776 -1378 956 -1366
rect -618 -1424 -244 -1420
rect 776 -1424 836 -1378
rect -618 -1442 836 -1424
rect 926 -1442 956 -1378
rect -618 -1444 956 -1442
rect -618 -1522 -572 -1444
rect -294 -1446 956 -1444
rect 1174 -1376 1334 -1366
rect 1174 -1440 1222 -1376
rect 1312 -1440 1334 -1376
rect 1174 -1446 1334 -1440
rect 2366 -1382 2480 -1372
rect 2366 -1442 2404 -1382
rect 2472 -1442 2480 -1382
rect 2366 -1444 2480 -1442
rect 2788 -1384 2852 -1374
rect -294 -1452 954 -1446
rect 1222 -1450 1312 -1446
rect 2404 -1452 2472 -1444
rect -294 -1522 -244 -1452
rect 2788 -1454 2852 -1444
rect -618 -1548 -244 -1522
rect 4718 -1712 4846 -1702
rect 6070 -1708 6444 -1696
rect 6070 -1710 6094 -1708
rect 6408 -1710 6444 -1708
rect 6070 -1770 6092 -1710
rect 6410 -1712 6444 -1710
rect 6434 -1770 6444 -1712
rect 6070 -1780 6444 -1770
rect 4718 -1800 4846 -1790
rect -144 -1936 6022 -1926
rect -144 -2124 6022 -2114
<< via2 >>
rect -232 1330 5994 1534
rect 2446 828 2508 884
rect -636 398 -374 458
rect -1470 -984 -1466 -858
rect -1466 -984 -1412 -858
rect -608 160 -328 238
rect 2434 192 2508 252
rect 2822 190 2892 248
rect 4746 -156 4874 -80
rect 6090 -144 6428 -88
rect 2764 -798 2872 -732
rect -440 -1232 -224 -1176
rect -572 -1522 -294 -1444
rect 2404 -1386 2472 -1382
rect 2404 -1438 2472 -1386
rect 2788 -1390 2852 -1384
rect 2788 -1444 2852 -1390
rect 4718 -1790 4846 -1712
rect 6092 -1712 6094 -1710
rect 6094 -1712 6408 -1710
rect 6408 -1712 6410 -1710
rect 6092 -1770 6434 -1712
rect -144 -2114 6022 -1936
<< metal3 >>
rect -242 1294 -232 1576
rect 6000 1294 6010 1576
rect 2438 894 2524 896
rect 2430 884 2524 894
rect 2430 866 2446 884
rect 2428 828 2446 866
rect 2508 828 2524 884
rect 2428 824 2524 828
rect 2428 778 2518 824
rect -476 738 -466 744
rect -500 658 -466 738
rect -476 644 -466 658
rect -366 738 -356 744
rect 2428 738 2508 778
rect -366 658 2508 738
rect -366 644 -356 658
rect -660 460 -344 466
rect -660 458 2506 460
rect -660 398 -636 458
rect -374 398 2506 458
rect -660 388 2506 398
rect -660 384 -344 388
rect 2434 274 2506 388
rect 2410 252 2528 274
rect -642 238 -302 246
rect -642 221 -608 238
rect -1130 160 -608 221
rect -328 160 -302 238
rect 2410 192 2434 252
rect 2508 192 2528 252
rect 2410 184 2528 192
rect 2796 248 2914 274
rect 2796 190 2822 248
rect 2892 190 2914 248
rect 2796 184 2914 190
rect -1130 155 -302 160
rect -1480 -858 -1398 -838
rect -1480 -984 -1470 -858
rect -1412 -887 -1398 -858
rect -1130 -887 -1064 155
rect -642 140 -302 155
rect 2812 -80 2892 184
rect -1412 -953 -1064 -887
rect -631 -128 2892 -80
rect 4736 -80 4884 -75
rect -631 -158 2890 -128
rect 4736 -156 4746 -80
rect 4874 -82 4884 -80
rect 6068 -82 6448 -78
rect 4874 -88 6449 -82
rect 4874 -144 6090 -88
rect 6428 -144 6449 -88
rect 4874 -152 6449 -144
rect 4874 -156 4944 -152
rect 6068 -154 6448 -152
rect -1412 -984 -1398 -953
rect -1480 -1004 -1398 -984
rect -1472 -1732 -1412 -1004
rect -631 -1420 -553 -158
rect 4736 -161 4884 -156
rect 2754 -732 2882 -727
rect 2754 -798 2764 -732
rect 2872 -798 2882 -732
rect 2754 -803 2882 -798
rect -470 -988 -460 -890
rect -354 -908 -344 -890
rect 2790 -908 2850 -803
rect -354 -968 2850 -908
rect -354 -988 -344 -968
rect -478 -1173 -190 -1162
rect -478 -1176 2462 -1173
rect -478 -1232 -440 -1176
rect -224 -1232 2462 -1176
rect -478 -1235 2462 -1232
rect -478 -1246 -190 -1235
rect 2400 -1356 2462 -1235
rect 2366 -1382 2482 -1356
rect 2798 -1358 2858 -1356
rect -631 -1444 -244 -1420
rect 2366 -1438 2404 -1382
rect 2472 -1438 2482 -1382
rect 2366 -1444 2482 -1438
rect 2772 -1384 2886 -1358
rect 2772 -1444 2788 -1384
rect 2852 -1444 2886 -1384
rect -631 -1522 -572 -1444
rect -294 -1522 -244 -1444
rect 2772 -1450 2886 -1444
rect -631 -1541 -244 -1522
rect -618 -1548 -244 -1541
rect 2798 -1732 2858 -1450
rect -1472 -1792 2858 -1732
rect 4708 -1712 4856 -1707
rect 6070 -1710 6444 -1696
rect 6070 -1712 6092 -1710
rect 6410 -1712 6444 -1710
rect 4708 -1790 4718 -1712
rect 4846 -1770 6092 -1712
rect 6434 -1770 6444 -1712
rect 4846 -1780 6444 -1770
rect 4846 -1790 4856 -1780
rect 4708 -1795 4856 -1790
rect -154 -1931 6028 -1896
rect -154 -1936 6032 -1931
rect -154 -2114 -144 -1936
rect 6022 -2114 6032 -1936
rect -154 -2119 6032 -2114
<< via3 >>
rect -232 1534 6000 1576
rect -232 1330 5994 1534
rect 5994 1330 6000 1534
rect -232 1294 6000 1330
rect -466 644 -366 744
rect -460 -988 -354 -890
<< metal4 >>
rect -232 1577 6022 1614
rect -233 1576 6022 1577
rect -233 1556 -232 1576
rect -276 1318 -232 1556
rect -233 1294 -232 1318
rect 6000 1294 6022 1576
rect -233 1293 6022 1294
rect -232 1228 6022 1293
rect -232 1214 4944 1228
rect 5714 1214 6022 1228
rect -467 744 -365 745
rect -467 644 -466 744
rect -366 644 -365 744
rect -467 643 -365 644
rect -466 -790 -366 643
rect -466 -890 -352 -790
rect -466 -984 -460 -890
rect -461 -988 -460 -984
rect -354 -984 -352 -890
rect -354 -988 -353 -984
rect -461 -989 -353 -988
use comparator_full_compact  comparator_full_compact_0
timestamp 1698871213
transform 1 0 622 0 1 -292
box -794 -4 5299 1494
use comparator_full_compact  comparator_full_compact_1
timestamp 1698871213
transform 1 0 592 0 1 -1922
box -794 -4 5299 1494
use reference  reference_0
timestamp 1698913862
transform 1 0 -2500 0 1 -1085
box -32 -858 1956 500
use sky130_fd_pr__nfet_01v8_GWFSUW  sky130_fd_pr__nfet_01v8_GWFSUW_0
timestamp 1698873245
transform 1 0 389 0 1 -442
box -413 -130 413 130
use sky130_fd_pr__nfet_01v8_GWFSUW  sky130_fd_pr__nfet_01v8_GWFSUW_1
timestamp 1698873245
transform 1 0 1283 0 1 -446
box -413 -130 413 130
use sky130_fd_pr__nfet_01v8_GWFSUW  sky130_fd_pr__nfet_01v8_GWFSUW_2
timestamp 1698873245
transform 1 0 2241 0 1 -444
box -413 -130 413 130
use sky130_fd_pr__nfet_01v8_GWFSUW  sky130_fd_pr__nfet_01v8_GWFSUW_3
timestamp 1698873245
transform 1 0 3199 0 1 -444
box -413 -130 413 130
use sky130_fd_pr__nfet_01v8_GWFSUW  sky130_fd_pr__nfet_01v8_GWFSUW_4
timestamp 1698873245
transform 1 0 4181 0 1 -446
box -413 -130 413 130
use sky130_fd_pr__nfet_01v8_GWFSUW  sky130_fd_pr__nfet_01v8_GWFSUW_5
timestamp 1698873245
transform 1 0 5123 0 1 -446
box -413 -130 413 130
use xnor  xnor_0 ~/Desktop/charge_pumps2/layout_files2
timestamp 1698771789
transform 1 0 6348 0 1 -1100
box -162 -48 2166 592
<< labels >>
rlabel metal2 -258 -1435 -258 -1435 1 Vc-
rlabel metal2 -253 -1302 -253 -1302 1 V+
rlabel via2 -289 -1211 -289 -1211 1 V-
rlabel metal3 -373 430 -373 430 1 V-
rlabel metal2 -369 312 -369 312 1 V+
rlabel via2 -380 200 -380 200 1 Vc+
rlabel metal3 -358 -112 -358 -112 1 Vc-
rlabel via2 6269 -129 6269 -129 1 Q2
rlabel via2 6329 -1756 6329 -1756 1 Q
rlabel metal1 -1384 428 -1384 428 1 V-
rlabel metal2 -692 -1088 -692 -1088 1 V+
port 5 n
rlabel metal1 6088 -566 6088 -566 1 q2
port 6 n
rlabel metal1 6088 -1304 6088 -1304 1 q
port 7 n
rlabel metal1 8530 -782 8530 -782 1 enable
port 8 n
rlabel metal4 -418 -746 -418 -746 1 clk
port 9 n
rlabel space -1348 -1526 -1348 -1526 1 vref-
rlabel metal1 -736 -1574 -736 -1574 1 vref-
rlabel metal1 -1440 436 -1440 436 1 V-
port 10 n
<< end >>
