magic
tech sky130A
magscale 1 2
timestamp 1698871213
<< locali >>
rect -3086 3526 -3000 3662
rect -1934 3528 -1848 3664
rect -1424 3620 -1218 3774
rect -900 3772 -712 3776
rect -1418 3494 -1230 3496
rect -3258 3380 -3100 3470
rect -2990 3386 -2832 3476
rect -2094 3386 -1952 3464
rect -1824 3388 -1682 3466
rect -916 3342 -710 3496
rect -3290 3196 -3158 3232
rect -2930 3196 -1678 3232
rect -3290 3166 -1678 3196
<< viali >>
rect -3158 3196 -2930 3232
rect -3174 2864 -3060 2974
rect -438 1032 -370 3064
<< metal1 >>
rect -1172 4012 -1162 4112
rect -1088 4012 -1078 4112
rect -3035 3966 -2781 3975
rect -3036 3936 -2781 3966
rect -3036 3664 -2992 3936
rect -3036 3620 -2148 3664
rect -2330 3562 -2320 3586
rect -2690 3522 -2320 3562
rect -2234 3522 -2224 3586
rect -2584 3474 -2538 3486
rect -2192 3478 -2148 3620
rect -1496 3538 -632 3582
rect -484 3538 -118 3582
rect -2612 3386 -2602 3474
rect -2540 3386 -2530 3474
rect -3170 3236 -2918 3238
rect -3293 3232 -2918 3236
rect -3293 3196 -3158 3232
rect -2930 3196 -2918 3232
rect -3293 3161 -2918 3196
rect -3202 2974 -3036 3161
rect -2716 3064 -2656 3342
rect -2584 3167 -2538 3386
rect -2194 3247 -2148 3478
rect -2194 3201 763 3247
rect -2584 3121 775 3167
rect -444 3064 -364 3076
rect -2716 3004 -438 3064
rect -3202 2864 -3174 2974
rect -3060 2864 -3036 2974
rect -3202 2842 -3036 2864
rect -448 1032 -438 3004
rect -370 1032 -360 3064
rect -444 1020 -364 1032
<< via1 >>
rect -1162 4012 -1088 4112
rect -2320 3522 -2234 3586
rect -2602 3386 -2540 3474
rect -3174 2864 -3060 2974
rect -438 1032 -370 3064
<< metal2 >>
rect -2180 3912 -2144 4186
rect -1162 4112 -1088 4122
rect -1162 4002 -1088 4012
rect -2602 3876 -2144 3912
rect -2602 3484 -2566 3876
rect -1121 3811 -1091 4002
rect -2304 3781 -1091 3811
rect -2304 3596 -2274 3781
rect -2320 3586 -2234 3596
rect -2320 3512 -2234 3522
rect -2602 3474 -2540 3484
rect -2602 3376 -2540 3386
rect -438 3064 -370 3074
rect -3174 2974 -3060 2984
rect -3174 2854 -3060 2864
rect -438 1022 -370 1032
<< via2 >>
rect -3174 2864 -3060 2974
rect -438 1032 -370 3064
<< metal3 >>
rect -448 3064 -360 3069
rect -3202 2844 -3192 2988
rect -3046 2844 -3036 2988
rect -448 1032 -438 3064
rect -370 1032 -360 3064
rect -448 1027 -360 1032
<< via3 >>
rect -3192 2974 -3046 2988
rect -3192 2864 -3174 2974
rect -3174 2864 -3060 2974
rect -3060 2864 -3046 2974
rect -3192 2844 -3046 2864
<< metal4 >>
rect -3202 2988 -3036 3230
rect -3202 2844 -3192 2988
rect -3046 2844 -2462 2988
rect -3202 2842 -3036 2844
use cmfb  cmfb_0
timestamp 1698789667
transform 1 0 -3134 0 1 2875
box 203 439 3639 2056
use sky130_fd_pr__nfet_01v8_53744R  sky130_fd_pr__nfet_01v8_53744R_0
timestamp 1698787694
transform 0 1 -809 -1 0 3560
box -246 -310 246 310
use sky130_fd_pr__nfet_01v8_53744R  sky130_fd_pr__nfet_01v8_53744R_1
timestamp 1698787694
transform 0 1 -1323 -1 0 3560
box -246 -310 246 310
use sky130_fd_pr__pfet_01v8_TM5SY6  sky130_fd_pr__pfet_01v8_TM5SY6_0
timestamp 1698155087
transform 1 0 -2275 0 1 3430
box -246 -269 246 269
use sky130_fd_pr__pfet_01v8_TM5SY6  sky130_fd_pr__pfet_01v8_TM5SY6_1
timestamp 1698155087
transform 1 0 -2661 0 1 3430
box -246 -269 246 269
use sky130_fd_pr__pfet_01v8_TM5SY6  sky130_fd_pr__pfet_01v8_TM5SY6_2
timestamp 1698155087
transform 1 0 -3047 0 1 3430
box -246 -269 246 269
use sky130_fd_pr__pfet_01v8_TM5SY6  sky130_fd_pr__pfet_01v8_TM5SY6_3
timestamp 1698155087
transform 1 0 -1889 0 1 3430
box -246 -269 246 269
use sky130_fd_pr__cap_mim_m3_1_4PHTN9  XC3
timestamp 1697610037
transform 1 0 -1539 0 1 2044
box -1186 -1040 1186 1040
<< end >>
