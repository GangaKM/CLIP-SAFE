magic
tech sky130A
magscale 1 2
timestamp 1698765726
<< nwell >>
rect -3654 2366 -2708 2420
rect -3654 1456 -2696 2366
rect -3654 568 -2708 1456
rect -3312 542 -3024 568
rect -3018 556 -2720 568
rect -396 566 184 2640
rect -1728 302 -1042 488
rect -2748 12 -1042 302
rect -1728 10 -1042 12
<< pwell >>
rect -3176 3480 -3114 4296
<< psubdiff >>
rect 426 3536 564 3564
rect 426 3468 460 3536
rect 524 3468 564 3536
rect 426 3440 564 3468
<< nsubdiff >>
rect -18 2512 104 2540
rect -18 2466 10 2512
rect 72 2466 104 2512
rect -18 2430 104 2466
rect -3618 1312 -3498 1338
rect -3618 1250 -3594 1312
rect -3528 1250 -3498 1312
rect -3618 1226 -3498 1250
rect -1502 404 -1394 430
rect -1502 360 -1480 404
rect -1428 360 -1394 404
rect -1502 332 -1394 360
<< psubdiffcont >>
rect 460 3468 524 3536
<< nsubdiffcont >>
rect 10 2466 72 2512
rect -3594 1250 -3528 1312
rect -1480 360 -1428 404
<< poly >>
rect 920 3008 950 3036
rect 822 2970 950 3008
rect 3686 2710 3716 2746
rect 3612 2680 3716 2710
rect -3274 1246 -3244 1346
rect -3274 1216 -3208 1246
rect -2800 944 -2720 946
rect -2800 916 -2716 944
rect -2752 816 -2716 916
rect -362 692 -330 790
rect -362 662 -300 692
<< locali >>
rect 444 3536 560 3558
rect 444 3468 458 3536
rect 524 3468 560 3536
rect 444 3448 560 3468
rect -2908 2916 -2766 2998
rect -2524 2918 -2382 3000
rect 3421 2814 3471 2915
rect 3421 2764 3576 2814
rect -18 2512 104 2540
rect -18 2466 10 2512
rect 72 2466 104 2512
rect -18 2430 104 2466
rect -3618 1312 -3498 1338
rect -3618 1250 -3594 1312
rect -3528 1250 -3498 1312
rect -3618 1226 -3498 1250
rect -1502 404 -1394 430
rect -1502 360 -1480 404
rect -1428 360 -1394 404
rect -1502 332 -1394 360
<< viali >>
rect -3802 4536 4658 4752
rect 458 3468 460 3536
rect 460 3468 524 3536
rect -1684 2750 782 2796
rect 10 2466 72 2512
rect -3594 1250 -3528 1312
rect -1478 360 -1428 404
rect -3800 -454 4732 -178
<< metal1 >>
rect -3835 4752 4779 4979
rect -3835 4536 -3802 4752
rect 4658 4536 4779 4752
rect -3835 4427 4779 4536
rect -3410 4404 640 4427
rect -3410 2770 -3346 4404
rect -3264 4326 -3224 4404
rect -3266 3706 -3224 4326
rect -3266 3702 -3226 3706
rect -3186 3554 -3176 4370
rect -3114 3554 -3104 4370
rect -3068 4323 -3028 4404
rect -3068 3608 -3024 4323
rect 312 4312 640 4404
rect 452 3536 530 3548
rect 38 3452 48 3506
rect 152 3452 162 3506
rect 452 3468 458 3536
rect 524 3468 530 3536
rect 452 3456 530 3468
rect 458 3408 524 3456
rect 3588 3442 3598 3500
rect 3704 3442 3714 3500
rect 3867 3470 4507 3507
rect -946 3160 -936 3216
rect -754 3186 -744 3216
rect -754 3160 -672 3186
rect -780 3112 -672 3160
rect 6 3114 36 3340
rect 232 3258 712 3408
rect 382 3246 680 3258
rect 132 3156 958 3204
rect 1076 3118 1208 3176
rect 1086 3116 1208 3118
rect -786 3084 -680 3096
rect -786 3068 -682 3084
rect 2 3054 998 3114
rect 1086 3086 1174 3116
rect 1086 3040 1148 3086
rect -1466 2972 -1456 3028
rect -1274 2972 -1264 3028
rect 50 2968 876 3016
rect 810 2932 852 2968
rect 1086 2932 1146 3040
rect -14 2872 1146 2932
rect 3618 2872 4128 2908
rect 3618 2868 3890 2872
rect -1684 2802 794 2822
rect -3410 2690 -3300 2770
rect -1696 2750 -1684 2802
rect 784 2750 794 2802
rect 3542 2762 3960 2824
rect -1696 2744 794 2750
rect -1696 2730 772 2744
rect -3606 1312 -3516 1318
rect -3410 1312 -3346 2690
rect -2630 2689 -1692 2702
rect -2755 2572 -2702 2679
rect -2640 2629 -2630 2689
rect -2002 2629 -1692 2689
rect 523 2653 1887 2699
rect 3516 2656 3786 2706
rect -650 2542 -556 2590
rect -362 2530 -330 2592
rect -204 2566 68 2568
rect -3296 2246 -3256 2328
rect -3296 2194 -3252 2246
rect -3606 1250 -3594 1312
rect -3528 1250 -3346 1312
rect -3292 1618 -3252 2194
rect -3292 1348 -3264 1618
rect -3292 1304 -3244 1348
rect -3606 1244 -3516 1250
rect -3410 496 -3346 1250
rect -3284 720 -3244 1304
rect -3182 730 -3124 2292
rect -3074 2142 -2934 2344
rect -3084 1514 -2934 2142
rect -3194 584 -3124 730
rect -3074 634 -2934 1514
rect -3072 622 -3032 634
rect -3194 496 -3128 584
rect -2870 496 -2812 2344
rect -366 2302 -328 2530
rect -479 2249 -406 2299
rect -372 2244 -322 2302
rect -2760 2202 -2708 2210
rect -2768 796 -2758 2202
rect -2694 796 -2684 2202
rect -372 2138 -321 2244
rect -371 2083 -321 2138
rect -270 2148 -212 2566
rect -204 2534 78 2566
rect -22 2518 78 2534
rect -22 2512 84 2518
rect -22 2466 10 2512
rect 72 2466 84 2512
rect -22 2462 84 2466
rect -2 2460 84 2462
rect 1841 2461 1887 2653
rect 2158 2470 2168 2536
rect 2262 2470 2272 2536
rect -152 2324 -112 2434
rect -476 1508 -400 1556
rect -366 750 -324 2083
rect -270 2010 -216 2148
rect -160 2028 -110 2324
rect -366 746 -328 750
rect -270 612 -206 2010
rect -152 700 -112 2028
rect -152 656 54 700
rect -260 496 -206 612
rect -3924 404 -112 496
rect -3924 360 -1478 404
rect -1428 360 -112 404
rect -3924 346 -112 360
rect -3924 340 -2354 346
rect -1338 340 -112 346
rect -3412 295 -3344 340
rect -3845 257 -2947 295
rect -2803 294 -2371 295
rect -3845 84 -3807 257
rect -3590 240 -2948 257
rect -2803 246 -1128 294
rect -2803 245 -2371 246
rect -3728 130 -2922 194
rect -3690 84 -3048 94
rect -3845 46 -3048 84
rect -3690 44 -3048 46
rect -2964 -56 -2926 130
rect -2803 104 -2753 245
rect -1100 192 -1062 340
rect -1028 338 -112 340
rect -724 273 -676 338
rect -1130 186 -1062 192
rect -2694 130 -1062 186
rect -975 223 -107 273
rect -2694 126 -1066 130
rect -2806 66 -2753 104
rect -975 72 -925 223
rect -94 176 -56 190
rect -872 126 -52 176
rect -2666 66 -1342 70
rect -2806 22 -1342 66
rect -975 22 -186 72
rect -2806 16 -2624 22
rect -2806 -56 -2754 16
rect -1420 -56 -1382 -54
rect -94 -56 -56 126
rect 10 -56 54 656
rect 1818 -56 2110 2182
rect -3834 -172 4728 -56
rect -3834 -178 4744 -172
rect -3834 -454 -3800 -178
rect 4732 -454 4744 -178
rect -3834 -460 4744 -454
rect -3834 -570 4728 -460
<< via1 >>
rect -3802 4536 4658 4752
rect -3176 3554 -3114 4370
rect 48 3452 152 3506
rect 3598 3442 3704 3500
rect -936 3160 -754 3216
rect -1456 2972 -1274 3028
rect -1684 2796 784 2802
rect -1684 2750 782 2796
rect 782 2750 784 2796
rect -2630 2629 -2002 2689
rect -2758 796 -2694 2202
rect 2168 2470 2262 2536
rect -3800 -454 4732 -178
<< metal2 >>
rect -3835 4752 4779 4979
rect -3835 4536 -3802 4752
rect 4658 4536 4779 4752
rect -3835 4427 4779 4536
rect -3176 4370 -3114 4380
rect -3176 3423 -3114 3554
rect 48 3506 152 3516
rect 48 3442 52 3452
rect 142 3442 152 3452
rect 3598 3500 3704 3510
rect 52 3430 142 3440
rect 3598 3432 3704 3442
rect -3176 3361 -2815 3423
rect -936 3216 -754 3226
rect -936 3150 -754 3160
rect -1456 3028 -1274 3038
rect -1456 2962 -1274 2972
rect -1684 2808 784 2818
rect -3564 2750 -1684 2808
rect -3564 2748 784 2750
rect -1684 2740 784 2748
rect -2630 2691 -2002 2699
rect -3583 2689 -2002 2691
rect -3583 2629 -2630 2689
rect -3583 2621 -2002 2629
rect -2630 2619 -2002 2621
rect 2158 2546 2250 2556
rect 2250 2536 2262 2546
rect 2250 2468 2262 2470
rect 2158 2460 2262 2468
rect 2158 2458 2250 2460
rect -2758 2210 -2694 2212
rect -2768 2202 -2694 2210
rect -2768 796 -2758 2202
rect 4256 1738 4712 1826
rect -2768 786 -2694 796
rect -2768 -56 -2698 786
rect -3800 -168 4728 -56
rect -3800 -178 4732 -168
rect -3800 -464 4732 -454
rect -3800 -570 4728 -464
<< via2 >>
rect -3802 4536 4658 4752
rect 52 3452 142 3506
rect 52 3440 142 3452
rect 3598 3442 3704 3500
rect -936 3160 -754 3216
rect -1456 2972 -1274 3028
rect -1684 2802 784 2808
rect -1684 2750 784 2802
rect 2158 2536 2250 2546
rect 2158 2470 2168 2536
rect 2168 2470 2250 2536
rect 2158 2468 2250 2470
rect -3800 -454 4732 -178
<< metal3 >>
rect -3835 4766 4779 4979
rect -3835 4494 -3802 4766
rect 4654 4752 4779 4766
rect 4658 4536 4779 4752
rect 4654 4494 4779 4536
rect -3835 4427 4779 4494
rect 32 3508 174 3512
rect -3555 3506 356 3508
rect -3555 3440 52 3506
rect 142 3440 356 3506
rect -3555 3434 356 3440
rect 3154 3500 3715 3508
rect 3154 3442 3598 3500
rect 3704 3442 3715 3500
rect 3154 3434 3715 3442
rect -960 3223 -780 3224
rect -3569 3216 -743 3223
rect -3569 3160 -936 3216
rect -754 3160 -743 3216
rect -3569 3154 -743 3160
rect -1466 3028 -1264 3033
rect -1466 3024 -1456 3028
rect -3558 2972 -1456 3024
rect -1274 2972 -1264 3028
rect -3558 2967 -1264 2972
rect -3558 2961 -1330 2967
rect -1510 2956 -1330 2961
rect -1684 2813 794 2822
rect -1694 2808 794 2813
rect -1694 2800 -1684 2808
rect -1726 2750 -1684 2800
rect 784 2750 794 2808
rect -1726 2745 794 2750
rect -1726 2732 768 2745
rect 700 2534 768 2732
rect 2148 2546 2260 2551
rect 2148 2534 2158 2546
rect 700 2468 2158 2534
rect 2250 2468 2260 2546
rect 700 2466 2260 2468
rect 2148 2463 2260 2466
rect 809 2182 4669 2257
rect -3834 -173 -3732 -56
rect -3834 -178 4742 -173
rect -3834 -454 -3800 -178
rect 4732 -454 4742 -178
rect -3834 -459 4742 -454
rect -3834 -570 -3732 -459
<< via3 >>
rect -3802 4752 4654 4766
rect -3802 4536 4658 4752
rect -3802 4494 4654 4536
rect -3800 -454 4732 -178
<< metal4 >>
rect -3835 4766 4779 4979
rect -3835 4494 -3802 4766
rect 4654 4752 4779 4766
rect 4658 4536 4779 4752
rect 4654 4494 4779 4536
rect -3835 4427 4779 4494
rect -3834 -177 -3732 -56
rect -3834 -178 4733 -177
rect -3834 -454 -3800 -178
rect 4732 -454 4733 -178
rect -3834 -455 4733 -454
rect -3834 -570 -3732 -455
<< via4 >>
rect -3800 -454 4732 -178
<< metal5 >>
rect -3834 -154 4728 -56
rect -3834 -178 4756 -154
rect -3834 -454 -3800 -178
rect 4732 -454 4756 -178
rect -3834 -478 4756 -454
rect -3834 -570 4728 -478
use firststage_compact  firststage_compact_0 ~/layout_files/differential_amplifier
timestamp 1698651669
transform 1 0 -43 0 1 -468
box -3293 1004 775 4931
use integrator_full_new_compact  integrator_full_new_compact_0 ~/layout_files/differential_amplifier
timestamp 1698651669
transform 1 0 386 0 1 3329
box -386 -3329 4003 1133
use sky130_fd_pr__nfet_01v8_647BNN  sky130_fd_pr__nfet_01v8_647BNN_0 ~/layout_files/differential_amplifier
timestamp 1698611618
transform 1 0 3749 0 1 2794
box -221 -130 221 130
use sky130_fd_pr__nfet_01v8_FU3CJE  sky130_fd_pr__nfet_01v8_FU3CJE_0 ~/layout_files/differential_amplifier
timestamp 1698611618
transform 1 0 503 0 1 3086
box -509 -130 509 130
use sky130_fd_pr__nfet_01v8_GWAZJ9  sky130_fd_pr__nfet_01v8_GWAZJ9_0 ~/layout_files/differential_amplifier
timestamp 1698611618
transform 1 0 -3323 0 1 164
box -413 -130 413 130
use sky130_fd_pr__nfet_01v8_GWAZJ9  sky130_fd_pr__nfet_01v8_GWAZJ9_1
timestamp 1698611618
transform 1 0 -469 0 1 152
box -413 -130 413 130
use sky130_fd_pr__nfet_01v8_GWXQMW  sky130_fd_pr__nfet_01v8_GWXQMW_0 ~/layout_files/differential_amplifier
timestamp 1698611618
transform 0 -1 -3146 1 0 3969
box -413 -130 413 130
use sky130_fd_pr__pfet_01v8_ACB9FB  sky130_fd_pr__pfet_01v8_ACB9FB_0 ~/layout_files/differential_amplifier
timestamp 1698611618
transform 0 -1 -3156 1 0 991
box -449 -142 449 142
use sky130_fd_pr__pfet_01v8_ACB9FB  sky130_fd_pr__pfet_01v8_ACB9FB_1
timestamp 1698611618
transform 0 -1 -3166 1 0 1883
box -449 -142 449 142
use sky130_fd_pr__pfet_01v8_ACB9FB  sky130_fd_pr__pfet_01v8_ACB9FB_2
timestamp 1698611618
transform 0 -1 -2840 1 0 1171
box -449 -142 449 142
use sky130_fd_pr__pfet_01v8_ACB9FB  sky130_fd_pr__pfet_01v8_ACB9FB_3
timestamp 1698611618
transform 0 -1 -2840 1 0 1939
box -449 -142 449 142
use sky130_fd_pr__pfet_01v8_DCBZKP  sky130_fd_pr__pfet_01v8_DCBZKP_0 ~/layout_files/differential_amplifier
timestamp 1698611618
transform 1 0 -1896 0 1 158
box -848 -142 848 142
use sky130_fd_pr__pfet_01v8_WMSBVE  sky130_fd_pr__pfet_01v8_WMSBVE_0 ~/layout_files/differential_amplifier
timestamp 1698611618
transform 0 -1 -240 1 0 1589
box -1025 -142 1025 142
<< labels >>
rlabel metal4 -3652 4448 -3652 4448 1 Vdd
rlabel metal5 -3228 -518 -3228 -518 1 gnd
rlabel metal1 -598 2574 -598 2574 1 Vbp
rlabel metal3 -3509 3189 -3509 3189 1 Vbias
rlabel metal3 -3509 2980 -3509 2980 1 Vs
rlabel metal2 -3490 2771 -3490 2771 1 vd2
rlabel metal2 -3506 2656 -3506 2656 1 vd1
rlabel metal1 4425 3485 4425 3485 1 Vcmref
rlabel metal2 4641 1770 4641 1770 1 vo1
rlabel metal3 4575 2201 4575 2201 1 vo2
rlabel metal3 -3510 3452 -3510 3452 1 Vcm_ref
<< end >>
