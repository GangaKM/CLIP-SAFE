magic
tech sky130A
magscale 1 2
timestamp 1698762467
<< error_p >>
rect 132733 85585 132747 85607
rect 132761 85606 132775 85607
rect 132733 83499 132747 83521
rect 132761 83520 132775 83521
rect 132731 81405 132745 81427
rect 132759 81426 132773 81427
rect 132731 79323 132745 79345
rect 132759 79344 132773 79345
rect 132731 77225 132745 77247
rect 132759 77246 132773 77247
rect 132805 75135 132819 75157
rect 132833 75156 132847 75157
rect 132807 73041 132821 73063
rect 132835 73062 132849 73063
rect 132485 -73241 132499 -73219
rect 132513 -73241 132527 -73240
rect 132483 -75335 132497 -75313
rect 132511 -75335 132525 -75334
rect 132409 -77425 132423 -77403
rect 132437 -77425 132451 -77424
rect 132409 -79523 132423 -79501
rect 132437 -79523 132451 -79522
rect 132409 -81605 132423 -81583
rect 132437 -81605 132451 -81604
rect 132411 -83699 132425 -83677
rect 132439 -83699 132453 -83698
rect 132411 -85785 132425 -85763
rect 132439 -85785 132453 -85784
<< metal1 >>
rect -1034 41744 -474 41752
rect -1034 41716 308 41744
rect -1034 -41894 -474 41716
rect -352 -41290 208 41136
rect -1034 -41922 50 -41894
rect -1034 -41926 -474 -41922
use comparator_final_compact  comparator_final_compact_0 ~/layout_files/differential_amplifier
timestamp 1698761357
transform -1 0 8823 0 1 -19510
box -2566 -2214 8653 1614
use reconfigurable_CP  reconfigurable_CP_0
timestamp 1698762467
transform 1 0 16242 0 -1 63194
box -16084 -36096 128734 63194
use reconfigurable_CP  reconfigurable_CP_1
timestamp 1698762467
transform 1 0 15920 0 1 -63372
box -16084 -36096 128734 63194
<< end >>
