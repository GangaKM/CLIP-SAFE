* SPICE3 file created from reconfigurable_CP.ext - technology: sky130A

.subckt sky130_fd_pr__cap_mim_m3_1_MH6KF8 c1_n1046_n900# m3_n1086_n940# VSUBS
X0 c1_n1046_n900# m3_n1086_n940# sky130_fd_pr__cap_mim_m3_1 l=9 w=9
C0 m3_n1086_n940# c1_n1046_n900# 7.78f
C1 m3_n1086_n940# VSUBS 3.31f
.ends

.subckt sky130_fd_pr__pfet_01v8_FXZ64Q a_n73_n126# w_n109_n188# a_15_n126# a_n15_n152#
+ VSUBS
X0 a_15_n126# a_n15_n152# a_n73_n126# w_n109_n188# sky130_fd_pr__pfet_01v8 ad=0.365 pd=3.1 as=0.365 ps=3.1 w=1.26 l=0.15
.ends

.subckt sky130_fd_pr__nfet_01v8_DQBD8A a_15_n42# a_n15_n68# a_n73_n42# VSUBS
X0 a_15_n42# a_n15_n68# a_n73_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
.ends

.subckt buffer_digital m1_304_98# a_116_148# m1_n2_474# sky130_fd_pr__pfet_01v8_FXZ64Q_1/w_n109_n188#
+ a_n274_130# m1_n2_0# m1_216_0# VSUBS
Xsky130_fd_pr__pfet_01v8_FXZ64Q_0 m1_n2_474# sky130_fd_pr__pfet_01v8_FXZ64Q_1/w_n109_n188#
+ a_116_148# a_n274_130# VSUBS sky130_fd_pr__pfet_01v8_FXZ64Q
Xsky130_fd_pr__pfet_01v8_FXZ64Q_1 m1_n2_474# sky130_fd_pr__pfet_01v8_FXZ64Q_1/w_n109_n188#
+ m1_304_98# a_116_148# VSUBS sky130_fd_pr__pfet_01v8_FXZ64Q
Xsky130_fd_pr__nfet_01v8_DQBD8A_0 a_116_148# a_n274_130# m1_n2_0# VSUBS sky130_fd_pr__nfet_01v8_DQBD8A
Xsky130_fd_pr__nfet_01v8_DQBD8A_1 m1_304_98# a_116_148# m1_216_0# VSUBS sky130_fd_pr__nfet_01v8_DQBD8A
.ends

.subckt sky130_fd_pr__nfet_01v8_D4CMYK a_15_n130# a_63_n42# a_n177_n130# a_255_n42#
+ a_n129_n42# a_111_64# a_n321_n42# a_159_n42# a_n81_64# a_n273_64# a_351_n42# a_207_n130#
+ a_303_64# a_n33_n42# a_n369_n130# a_n225_n42# a_n413_n42# VSUBS
X0 a_63_n42# a_15_n130# a_n33_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X1 a_n33_n42# a_n81_64# a_n129_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X2 a_351_n42# a_303_64# a_255_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X3 a_159_n42# a_111_64# a_63_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X4 a_255_n42# a_207_n130# a_159_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X5 a_n321_n42# a_n369_n130# a_n413_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X6 a_n225_n42# a_n273_64# a_n321_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X7 a_n129_n42# a_n177_n130# a_n225_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
.ends

.subckt sky130_fd_pr__pfet_01v8_4ZKXAA a_63_n42# a_n417_n42# a_303_n139# w_n545_n142#
+ a_255_n42# a_n465_n139# a_n129_n42# a_111_n139# a_447_n42# a_n273_n139# a_n177_73#
+ a_n321_n42# a_207_73# a_n509_n42# a_159_n42# a_15_73# a_n81_n139# a_351_n42# a_n33_n42#
+ a_n369_73# a_n225_n42# a_399_73# VSUBS
X0 a_n33_n42# a_n81_n139# a_n129_n42# w_n545_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X1 a_351_n42# a_303_n139# a_255_n42# w_n545_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X2 a_159_n42# a_111_n139# a_63_n42# w_n545_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X3 a_255_n42# a_207_73# a_159_n42# w_n545_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X4 a_447_n42# a_399_73# a_351_n42# w_n545_n142# sky130_fd_pr__pfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X5 a_n321_n42# a_n369_73# a_n417_n42# w_n545_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X6 a_n225_n42# a_n273_n139# a_n321_n42# w_n545_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X7 a_n417_n42# a_n465_n139# a_n509_n42# w_n545_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X8 a_n129_n42# a_n177_73# a_n225_n42# w_n545_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X9 a_63_n42# a_15_73# a_n33_n42# w_n545_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
.ends

.subckt sky130_fd_pr__nfet_01v8_NJGC45 a_63_n42# a_15_64# a_n417_n42# a_111_n130#
+ a_n273_n130# a_255_n42# a_n129_n42# a_n369_64# a_399_64# a_447_n42# a_n81_n130#
+ a_n321_n42# a_n509_n42# a_159_n42# a_351_n42# a_n33_n42# a_303_n130# a_n225_n42#
+ a_n177_64# a_207_64# a_n465_n130# VSUBS
X0 a_63_n42# a_15_64# a_n33_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X1 a_n33_n42# a_n81_n130# a_n129_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X2 a_351_n42# a_303_n130# a_255_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X3 a_159_n42# a_111_n130# a_63_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X4 a_255_n42# a_207_64# a_159_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X5 a_447_n42# a_399_64# a_351_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X6 a_n321_n42# a_n369_64# a_n417_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X7 a_n417_n42# a_n465_n130# a_n509_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X8 a_n225_n42# a_n273_n130# a_n321_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X9 a_n129_n42# a_n177_64# a_n225_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
.ends

.subckt sky130_fd_pr__nfet_01v8_NJGLN5 a_n129_n130# a_n369_n42# a_1215_n130# a_543_64#
+ a_63_n130# a_159_64# a_n1089_n130# a_n849_n42# a_n417_64# a_n801_64# a_687_n42#
+ a_303_n42# a_1167_n42# a_n561_n42# a_n321_n130# a_n1041_n42# a_639_n130# a_n1185_64#
+ a_1023_n130# a_n1281_n130# a_n81_n42# a_399_n42# a_879_n42# a_n273_n42# a_735_64#
+ a_n753_n42# a_15_n42# a_n897_n130# a_n1233_n42# a_831_n130# a_447_n130# a_n609_64#
+ a_1071_n42# a_591_n42# a_1119_64# a_n993_64# a_207_n42# a_n465_n42# a_n945_n42#
+ a_351_64# a_783_n42# a_255_n130# a_n33_64# a_n225_64# a_n705_n130# a_1263_n42# a_927_64#
+ a_n177_n42# a_n657_n42# a_n1325_n42# a_n1137_n42# a_495_n42# a_111_n42# a_975_n42#
+ a_n513_n130# VSUBS
X0 a_303_n42# a_255_n130# a_207_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X1 a_591_n42# a_543_64# a_495_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X2 a_207_n42# a_159_64# a_111_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X3 a_399_n42# a_351_64# a_303_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X4 a_495_n42# a_447_n130# a_399_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X5 a_687_n42# a_639_n130# a_591_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X6 a_783_n42# a_735_64# a_687_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X7 a_975_n42# a_927_64# a_879_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X8 a_n1041_n42# a_n1089_n130# a_n1137_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X9 a_879_n42# a_831_n130# a_783_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X10 a_n1233_n42# a_n1281_n130# a_n1325_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X11 a_n1137_n42# a_n1185_64# a_n1233_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X12 a_n561_n42# a_n609_64# a_n657_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X13 a_1071_n42# a_1023_n130# a_975_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X14 a_1263_n42# a_1215_n130# a_1167_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X15 a_n945_n42# a_n993_64# a_n1041_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X16 a_n753_n42# a_n801_64# a_n849_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X17 a_n657_n42# a_n705_n130# a_n753_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X18 a_n465_n42# a_n513_n130# a_n561_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X19 a_n369_n42# a_n417_64# a_n465_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X20 a_1167_n42# a_1119_64# a_1071_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X21 a_n849_n42# a_n897_n130# a_n945_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X22 a_15_n42# a_n33_64# a_n81_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X23 a_111_n42# a_63_n130# a_15_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X24 a_n273_n42# a_n321_n130# a_n369_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X25 a_n81_n42# a_n129_n130# a_n177_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X26 a_n177_n42# a_n225_64# a_n273_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
.ends

.subckt sky130_fd_pr__pfet_01v8_VR4B8J a_1119_157# a_783_n126# a_n81_n126# a_n849_n126#
+ a_399_n126# a_n1041_n126# a_351_157# a_495_n126# a_n945_n126# a_n33_157# a_n129_n223#
+ a_n513_n223# a_1215_n223# a_63_n223# a_n1089_n223# a_n225_157# a_591_n126# a_n657_n126#
+ a_207_n126# a_543_157# a_n1325_n126# a_n369_n126# a_n753_n126# a_n321_n223# a_303_n126#
+ a_1023_n223# a_639_n223# a_n1281_n223# a_n417_157# a_n465_n126# a_1167_n126# a_735_157#
+ a_15_n126# a_n561_n126# a_n993_157# a_n177_n126# a_n897_n223# w_n1361_n226# a_1263_n126#
+ a_879_n126# a_111_n126# a_831_n223# a_n609_157# a_447_n223# a_n273_n126# a_n1137_n126#
+ a_975_n126# a_927_157# a_n1185_157# a_n1233_n126# a_n801_157# a_1071_n126# a_687_n126#
+ a_255_n223# a_n705_n223# a_159_157# VSUBS
X0 a_n273_n126# a_n321_n223# a_n369_n126# w_n1361_n226# sky130_fd_pr__pfet_01v8 ad=0.208 pd=1.59 as=0.208 ps=1.59 w=1.26 l=0.15
X1 a_n1233_n126# a_n1281_n223# a_n1325_n126# w_n1361_n226# sky130_fd_pr__pfet_01v8 ad=0.208 pd=1.59 as=0.391 ps=3.14 w=1.26 l=0.15
X2 a_591_n126# a_543_157# a_495_n126# w_n1361_n226# sky130_fd_pr__pfet_01v8 ad=0.208 pd=1.59 as=0.208 ps=1.59 w=1.26 l=0.15
X3 a_n849_n126# a_n897_n223# a_n945_n126# w_n1361_n226# sky130_fd_pr__pfet_01v8 ad=0.208 pd=1.59 as=0.208 ps=1.59 w=1.26 l=0.15
X4 a_207_n126# a_159_157# a_111_n126# w_n1361_n226# sky130_fd_pr__pfet_01v8 ad=0.208 pd=1.59 as=0.208 ps=1.59 w=1.26 l=0.15
X5 a_n177_n126# a_n225_157# a_n273_n126# w_n1361_n226# sky130_fd_pr__pfet_01v8 ad=0.208 pd=1.59 as=0.208 ps=1.59 w=1.26 l=0.15
X6 a_n1137_n126# a_n1185_157# a_n1233_n126# w_n1361_n226# sky130_fd_pr__pfet_01v8 ad=0.208 pd=1.59 as=0.208 ps=1.59 w=1.26 l=0.15
X7 a_495_n126# a_447_n223# a_399_n126# w_n1361_n226# sky130_fd_pr__pfet_01v8 ad=0.208 pd=1.59 as=0.208 ps=1.59 w=1.26 l=0.15
X8 a_n561_n126# a_n609_157# a_n657_n126# w_n1361_n226# sky130_fd_pr__pfet_01v8 ad=0.208 pd=1.59 as=0.208 ps=1.59 w=1.26 l=0.15
X9 a_111_n126# a_63_n223# a_15_n126# w_n1361_n226# sky130_fd_pr__pfet_01v8 ad=0.208 pd=1.59 as=0.208 ps=1.59 w=1.26 l=0.15
X10 a_783_n126# a_735_157# a_687_n126# w_n1361_n226# sky130_fd_pr__pfet_01v8 ad=0.208 pd=1.59 as=0.208 ps=1.59 w=1.26 l=0.15
X11 a_1071_n126# a_1023_n223# a_975_n126# w_n1361_n226# sky130_fd_pr__pfet_01v8 ad=0.208 pd=1.59 as=0.208 ps=1.59 w=1.26 l=0.15
X12 a_399_n126# a_351_157# a_303_n126# w_n1361_n226# sky130_fd_pr__pfet_01v8 ad=0.208 pd=1.59 as=0.208 ps=1.59 w=1.26 l=0.15
X13 a_n465_n126# a_n513_n223# a_n561_n126# w_n1361_n226# sky130_fd_pr__pfet_01v8 ad=0.208 pd=1.59 as=0.208 ps=1.59 w=1.26 l=0.15
X14 a_687_n126# a_639_n223# a_591_n126# w_n1361_n226# sky130_fd_pr__pfet_01v8 ad=0.208 pd=1.59 as=0.208 ps=1.59 w=1.26 l=0.15
X15 a_n753_n126# a_n801_157# a_n849_n126# w_n1361_n226# sky130_fd_pr__pfet_01v8 ad=0.208 pd=1.59 as=0.208 ps=1.59 w=1.26 l=0.15
X16 a_975_n126# a_927_157# a_879_n126# w_n1361_n226# sky130_fd_pr__pfet_01v8 ad=0.208 pd=1.59 as=0.208 ps=1.59 w=1.26 l=0.15
X17 a_n81_n126# a_n129_n223# a_n177_n126# w_n1361_n226# sky130_fd_pr__pfet_01v8 ad=0.208 pd=1.59 as=0.208 ps=1.59 w=1.26 l=0.15
X18 a_15_n126# a_n33_157# a_n81_n126# w_n1361_n226# sky130_fd_pr__pfet_01v8 ad=0.208 pd=1.59 as=0.208 ps=1.59 w=1.26 l=0.15
X19 a_1263_n126# a_1215_n223# a_1167_n126# w_n1361_n226# sky130_fd_pr__pfet_01v8 ad=0.391 pd=3.14 as=0.208 ps=1.59 w=1.26 l=0.15
X20 a_n1041_n126# a_n1089_n223# a_n1137_n126# w_n1361_n226# sky130_fd_pr__pfet_01v8 ad=0.208 pd=1.59 as=0.208 ps=1.59 w=1.26 l=0.15
X21 a_n369_n126# a_n417_157# a_n465_n126# w_n1361_n226# sky130_fd_pr__pfet_01v8 ad=0.208 pd=1.59 as=0.208 ps=1.59 w=1.26 l=0.15
X22 a_n657_n126# a_n705_n223# a_n753_n126# w_n1361_n226# sky130_fd_pr__pfet_01v8 ad=0.208 pd=1.59 as=0.208 ps=1.59 w=1.26 l=0.15
X23 a_879_n126# a_831_n223# a_783_n126# w_n1361_n226# sky130_fd_pr__pfet_01v8 ad=0.208 pd=1.59 as=0.208 ps=1.59 w=1.26 l=0.15
X24 a_n945_n126# a_n993_157# a_n1041_n126# w_n1361_n226# sky130_fd_pr__pfet_01v8 ad=0.208 pd=1.59 as=0.208 ps=1.59 w=1.26 l=0.15
X25 a_1167_n126# a_1119_157# a_1071_n126# w_n1361_n226# sky130_fd_pr__pfet_01v8 ad=0.208 pd=1.59 as=0.208 ps=1.59 w=1.26 l=0.15
X26 a_303_n126# a_255_n223# a_207_n126# w_n1361_n226# sky130_fd_pr__pfet_01v8 ad=0.208 pd=1.59 as=0.208 ps=1.59 w=1.26 l=0.15
C0 w_n1361_n226# VSUBS 3.67f
.ends

.subckt buffer m1_n1188_2032# a_1504_1398# m1_n1188_1271# m5_n1320_776# a_n1158_1778#
+ a_1504_1860# a_1596_1398# w_1358_2156# m4_n1330_2222# VSUBS
Xsky130_fd_pr__nfet_01v8_NJGLN5_1 a_n1158_1778# m1_n1188_1271# a_n1158_1778# a_n1158_1778#
+ a_n1158_1778# a_n1158_1778# a_n1158_1778# a_1436_1552# a_n1158_1778# a_n1158_1778#
+ a_1436_1552# a_1436_1552# m1_n1188_1271# m1_n1188_1271# a_n1158_1778# a_1436_1552#
+ a_n1158_1778# a_n1158_1778# a_n1158_1778# a_n1158_1778# a_1436_1552# m1_n1188_1271#
+ a_1436_1552# a_1436_1552# a_n1158_1778# m1_n1188_1271# m1_n1188_1271# a_n1158_1778#
+ a_1436_1552# a_n1158_1778# a_n1158_1778# a_n1158_1778# a_1436_1552# m1_n1188_1271#
+ a_n1158_1778# a_n1158_1778# m1_n1188_1271# a_1436_1552# m1_n1188_1271# a_n1158_1778#
+ m1_n1188_1271# a_n1158_1778# a_n1158_1778# a_n1158_1778# a_n1158_1778# a_1436_1552#
+ a_n1158_1778# m1_n1188_1271# a_1436_1552# m1_n1188_1271# m1_n1188_1271# a_1436_1552#
+ a_1436_1552# m1_n1188_1271# a_n1158_1778# VSUBS sky130_fd_pr__nfet_01v8_NJGLN5
Xsky130_fd_pr__pfet_01v8_VR4B8J_1 a_n1158_1778# m1_n1188_2032# a_1436_1552# a_1436_1552#
+ m1_n1188_2032# a_1436_1552# a_n1158_1778# a_1436_1552# m1_n1188_2032# a_n1158_1778#
+ a_n1158_1778# a_n1158_1778# a_n1158_1778# a_n1158_1778# a_n1158_1778# a_n1158_1778#
+ m1_n1188_2032# a_1436_1552# m1_n1188_2032# a_n1158_1778# m1_n1188_2032# m1_n1188_2032#
+ m1_n1188_2032# a_n1158_1778# a_1436_1552# a_n1158_1778# a_n1158_1778# a_n1158_1778#
+ a_n1158_1778# a_1436_1552# m1_n1188_2032# a_n1158_1778# m1_n1188_2032# m1_n1188_2032#
+ a_n1158_1778# m1_n1188_2032# a_n1158_1778# w_1358_2156# a_1436_1552# a_1436_1552#
+ a_1436_1552# a_n1158_1778# a_n1158_1778# a_n1158_1778# a_1436_1552# m1_n1188_2032#
+ m1_n1188_2032# a_n1158_1778# a_n1158_1778# a_1436_1552# a_n1158_1778# a_1436_1552#
+ a_1436_1552# a_n1158_1778# a_n1158_1778# a_n1158_1778# VSUBS sky130_fd_pr__pfet_01v8_VR4B8J
X0 a_1504_1398# a_1436_1552# a_1596_1398# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X1 a_1504_1860# a_1436_1552# a_1596_1398# w_1358_2156# sky130_fd_pr__pfet_01v8 ad=0.208 pd=1.59 as=0.208 ps=1.59 w=1.26 l=0.15
X2 a_1596_1398# a_1436_1552# a_1504_1398# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X3 a_1596_1398# a_1436_1552# a_1504_1860# w_1358_2156# sky130_fd_pr__pfet_01v8 ad=0.208 pd=1.59 as=0.208 ps=1.59 w=1.26 l=0.15
X4 a_1596_1398# a_1436_1552# a_1504_1860# w_1358_2156# sky130_fd_pr__pfet_01v8 ad=0.391 pd=3.14 as=0.208 ps=1.59 w=1.26 l=0.15
X5 a_1596_1398# a_1436_1552# a_1504_1860# w_1358_2156# sky130_fd_pr__pfet_01v8 ad=0.208 pd=1.59 as=0.391 ps=3.14 w=1.26 l=0.15
X6 a_1596_1398# a_1436_1552# a_1504_1398# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X7 a_1504_1860# a_1436_1552# a_1596_1398# w_1358_2156# sky130_fd_pr__pfet_01v8 ad=0.208 pd=1.59 as=0.208 ps=1.59 w=1.26 l=0.15
X8 a_1596_1398# a_1436_1552# a_1504_1398# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X9 a_1504_1398# a_1436_1552# a_1596_1398# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X10 a_1504_1860# a_1436_1552# a_1596_1398# w_1358_2156# sky130_fd_pr__pfet_01v8 ad=0.208 pd=1.59 as=0.208 ps=1.59 w=1.26 l=0.15
X11 a_1596_1398# a_1436_1552# a_1504_1860# w_1358_2156# sky130_fd_pr__pfet_01v8 ad=0.208 pd=1.59 as=0.208 ps=1.59 w=1.26 l=0.15
X12 a_1504_1398# a_1436_1552# a_1596_1398# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X13 a_1596_1398# a_1436_1552# a_1504_1398# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X14 a_1596_1398# a_1436_1552# a_1504_1860# w_1358_2156# sky130_fd_pr__pfet_01v8 ad=0.208 pd=1.59 as=0.208 ps=1.59 w=1.26 l=0.15
X15 a_1504_1860# a_1436_1552# a_1596_1398# w_1358_2156# sky130_fd_pr__pfet_01v8 ad=0.208 pd=1.59 as=0.208 ps=1.59 w=1.26 l=0.15
X16 a_1504_1860# a_1436_1552# a_1596_1398# w_1358_2156# sky130_fd_pr__pfet_01v8 ad=0.208 pd=1.59 as=0.208 ps=1.59 w=1.26 l=0.15
X17 a_1504_1398# a_1436_1552# a_1596_1398# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X18 a_1596_1398# a_1436_1552# a_1504_1398# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X19 a_1596_1398# a_1436_1552# a_1504_1860# w_1358_2156# sky130_fd_pr__pfet_01v8 ad=0.208 pd=1.59 as=0.208 ps=1.59 w=1.26 l=0.15
X20 a_1596_1398# a_1436_1552# a_1504_1860# w_1358_2156# sky130_fd_pr__pfet_01v8 ad=0.208 pd=1.59 as=0.208 ps=1.59 w=1.26 l=0.15
X21 a_1504_1398# a_1436_1552# a_1596_1398# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X22 a_1596_1398# a_1436_1552# a_1504_1398# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X23 a_1504_1860# a_1436_1552# a_1596_1398# w_1358_2156# sky130_fd_pr__pfet_01v8 ad=0.208 pd=1.59 as=0.208 ps=1.59 w=1.26 l=0.15
X24 a_1504_1398# a_1436_1552# a_1596_1398# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X25 a_1504_1398# a_1436_1552# a_1596_1398# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X26 a_1596_1398# a_1436_1552# a_1504_1860# w_1358_2156# sky130_fd_pr__pfet_01v8 ad=0.208 pd=1.59 as=0.208 ps=1.59 w=1.26 l=0.15
X27 a_1596_1398# a_1436_1552# a_1504_1398# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X28 a_1504_1398# a_1436_1552# a_1596_1398# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X29 a_1596_1398# a_1436_1552# a_1504_1860# w_1358_2156# sky130_fd_pr__pfet_01v8 ad=0.208 pd=1.59 as=0.208 ps=1.59 w=1.26 l=0.15
X30 a_1504_1398# a_1436_1552# a_1596_1398# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X31 a_1596_1398# a_1436_1552# a_1504_1860# w_1358_2156# sky130_fd_pr__pfet_01v8 ad=0.208 pd=1.59 as=0.208 ps=1.59 w=1.26 l=0.15
X32 a_1596_1398# a_1436_1552# a_1504_1398# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X33 a_1596_1398# a_1436_1552# a_1504_1398# VSUBS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X34 a_1504_1860# a_1436_1552# a_1596_1398# w_1358_2156# sky130_fd_pr__pfet_01v8 ad=0.208 pd=1.59 as=0.208 ps=1.59 w=1.26 l=0.15
X35 a_1596_1398# a_1436_1552# a_1504_1398# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X36 a_1504_1398# a_1436_1552# a_1596_1398# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X37 a_1504_1860# a_1436_1552# a_1596_1398# w_1358_2156# sky130_fd_pr__pfet_01v8 ad=0.208 pd=1.59 as=0.208 ps=1.59 w=1.26 l=0.15
X38 a_1596_1398# a_1436_1552# a_1504_1860# w_1358_2156# sky130_fd_pr__pfet_01v8 ad=0.208 pd=1.59 as=0.208 ps=1.59 w=1.26 l=0.15
X39 a_1504_1398# a_1436_1552# a_1596_1398# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X40 a_1596_1398# a_1436_1552# a_1504_1398# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X41 a_1596_1398# a_1436_1552# a_1504_1398# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X42 a_1504_1860# a_1436_1552# a_1596_1398# w_1358_2156# sky130_fd_pr__pfet_01v8 ad=0.208 pd=1.59 as=0.208 ps=1.59 w=1.26 l=0.15
X43 a_1504_1398# a_1436_1552# a_1596_1398# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X44 a_1596_1398# a_1436_1552# a_1504_1860# w_1358_2156# sky130_fd_pr__pfet_01v8 ad=0.208 pd=1.59 as=0.208 ps=1.59 w=1.26 l=0.15
X45 a_1504_1860# a_1436_1552# a_1596_1398# w_1358_2156# sky130_fd_pr__pfet_01v8 ad=0.208 pd=1.59 as=0.208 ps=1.59 w=1.26 l=0.15
X46 a_1504_1398# a_1436_1552# a_1596_1398# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X47 a_1596_1398# a_1436_1552# a_1504_1860# w_1358_2156# sky130_fd_pr__pfet_01v8 ad=0.208 pd=1.59 as=0.208 ps=1.59 w=1.26 l=0.15
X48 a_1504_1860# a_1436_1552# a_1596_1398# w_1358_2156# sky130_fd_pr__pfet_01v8 ad=0.208 pd=1.59 as=0.208 ps=1.59 w=1.26 l=0.15
X49 a_1504_1860# a_1436_1552# a_1596_1398# w_1358_2156# sky130_fd_pr__pfet_01v8 ad=0.208 pd=1.59 as=0.208 ps=1.59 w=1.26 l=0.15
X50 a_1596_1398# a_1436_1552# a_1504_1398# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X51 a_1596_1398# a_1436_1552# a_1504_1398# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X52 a_1596_1398# a_1436_1552# a_1504_1860# w_1358_2156# sky130_fd_pr__pfet_01v8 ad=0.208 pd=1.59 as=0.208 ps=1.59 w=1.26 l=0.15
X53 a_1504_1860# a_1436_1552# a_1596_1398# w_1358_2156# sky130_fd_pr__pfet_01v8 ad=0.208 pd=1.59 as=0.208 ps=1.59 w=1.26 l=0.15
C0 a_1436_1552# w_1358_2156# 2.61f
C1 a_1596_1398# a_1504_1398# 2.65f
C2 a_1504_1860# a_1596_1398# 6.79f
C3 a_1436_1552# a_1596_1398# 2.21f
C4 m5_n1320_776# VSUBS 2.52f
C5 a_n1158_1778# VSUBS 7.08f
C6 a_1436_1552# VSUBS 8.93f
C7 w_1358_2156# VSUBS 5.14f
.ends

.subckt sky130_fd_pr__pfet_01v8_X4L24Q a_n33_n126# w_n353_n226# a_n317_n126# a_n177_157#
+ a_159_n126# a_111_n223# a_n273_n223# a_255_n126# a_n129_n126# a_n81_n223# a_63_n126#
+ a_n225_n126# a_15_157# a_207_157# VSUBS
X0 a_159_n126# a_111_n223# a_63_n126# w_n353_n226# sky130_fd_pr__pfet_01v8 ad=0.208 pd=1.59 as=0.208 ps=1.59 w=1.26 l=0.15
X1 a_n225_n126# a_n273_n223# a_n317_n126# w_n353_n226# sky130_fd_pr__pfet_01v8 ad=0.208 pd=1.59 as=0.391 ps=3.14 w=1.26 l=0.15
X2 a_63_n126# a_15_157# a_n33_n126# w_n353_n226# sky130_fd_pr__pfet_01v8 ad=0.208 pd=1.59 as=0.208 ps=1.59 w=1.26 l=0.15
X3 a_n129_n126# a_n177_157# a_n225_n126# w_n353_n226# sky130_fd_pr__pfet_01v8 ad=0.208 pd=1.59 as=0.208 ps=1.59 w=1.26 l=0.15
X4 a_n33_n126# a_n81_n223# a_n129_n126# w_n353_n226# sky130_fd_pr__pfet_01v8 ad=0.208 pd=1.59 as=0.208 ps=1.59 w=1.26 l=0.15
X5 a_255_n126# a_207_157# a_159_n126# w_n353_n226# sky130_fd_pr__pfet_01v8 ad=0.391 pd=3.14 as=0.208 ps=1.59 w=1.26 l=0.15
.ends

.subckt sky130_fd_pr__nfet_01v8_XJUN3E a_63_n42# a_15_64# a_111_n130# a_n273_n130#
+ a_255_n42# a_n129_n42# a_n317_n42# a_n81_n130# a_159_n42# a_n33_n42# a_n225_n42#
+ a_n177_64# a_207_64# VSUBS
X0 a_63_n42# a_15_64# a_n33_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X1 a_n33_n42# a_n81_n130# a_n129_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X2 a_159_n42# a_111_n130# a_63_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X3 a_255_n42# a_207_64# a_159_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X4 a_n225_n42# a_n273_n130# a_n317_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X5 a_n129_n42# a_n177_64# a_n225_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
.ends

.subckt and_gate a_514_134# w_n260_286# sky130_fd_pr__pfet_01v8_X4L24Q_0/VSUBS a_n162_206#
+ m1_748_n50#
Xsky130_fd_pr__pfet_01v8_X4L24Q_0 w_n260_286# w_n260_286# m1_748_n50# a_n78_396# w_n260_286#
+ a_n78_396# a_n78_396# m1_748_n50# m1_748_n50# a_n78_396# m1_748_n50# w_n260_286#
+ a_n78_396# a_n78_396# sky130_fd_pr__pfet_01v8_X4L24Q_0/VSUBS sky130_fd_pr__pfet_01v8_X4L24Q
Xsky130_fd_pr__nfet_01v8_XJUN3E_0 m1_748_n50# a_n78_396# a_n78_396# a_n78_396# m1_748_n50#
+ m1_748_n50# m1_748_n50# a_n78_396# sky130_fd_pr__pfet_01v8_X4L24Q_0/VSUBS sky130_fd_pr__pfet_01v8_X4L24Q_0/VSUBS
+ sky130_fd_pr__pfet_01v8_X4L24Q_0/VSUBS a_n78_396# a_n78_396# sky130_fd_pr__pfet_01v8_X4L24Q_0/VSUBS
+ sky130_fd_pr__nfet_01v8_XJUN3E
X0 a_n78_396# a_n162_206# w_n260_286# w_n260_286# sky130_fd_pr__pfet_01v8 ad=0.208 pd=1.59 as=0.208 ps=1.59 w=1.26 l=0.15
X1 sky130_fd_pr__pfet_01v8_X4L24Q_0/VSUBS a_n162_206# a_n78_n64# sky130_fd_pr__pfet_01v8_X4L24Q_0/VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X2 w_n260_286# a_n162_206# a_n78_396# w_n260_286# sky130_fd_pr__pfet_01v8 ad=0.208 pd=1.59 as=0.208 ps=1.59 w=1.26 l=0.15
X3 w_n260_286# a_n162_206# a_n78_396# w_n260_286# sky130_fd_pr__pfet_01v8 ad=0.208 pd=1.59 as=0.208 ps=1.59 w=1.26 l=0.15
X4 a_n78_396# a_n162_206# w_n260_286# w_n260_286# sky130_fd_pr__pfet_01v8 ad=0.195 pd=1.57 as=0.208 ps=1.59 w=1.26 l=0.15
X5 a_n78_396# a_514_134# a_n78_n64# sky130_fd_pr__pfet_01v8_X4L24Q_0/VSUBS sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0651 ps=0.73 w=0.42 l=0.15
X6 a_n78_n64# a_n162_206# sky130_fd_pr__pfet_01v8_X4L24Q_0/VSUBS sky130_fd_pr__pfet_01v8_X4L24Q_0/VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X7 w_n260_286# a_514_134# a_n78_396# w_n260_286# sky130_fd_pr__pfet_01v8 ad=0.365 pd=3.1 as=0.195 ps=1.57 w=1.26 l=0.15
X8 a_n78_396# a_n162_206# w_n260_286# w_n260_286# sky130_fd_pr__pfet_01v8 ad=0.208 pd=1.59 as=0.208 ps=1.59 w=1.26 l=0.15
X9 sky130_fd_pr__pfet_01v8_X4L24Q_0/VSUBS a_n162_206# a_n78_n64# sky130_fd_pr__pfet_01v8_X4L24Q_0/VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X10 w_n260_286# a_n162_206# a_n78_396# w_n260_286# sky130_fd_pr__pfet_01v8 ad=0.208 pd=1.59 as=0.391 ps=3.14 w=1.26 l=0.15
X11 sky130_fd_pr__pfet_01v8_X4L24Q_0/VSUBS a_n162_206# a_n78_n64# sky130_fd_pr__pfet_01v8_X4L24Q_0/VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X12 a_n78_n64# a_n162_206# sky130_fd_pr__pfet_01v8_X4L24Q_0/VSUBS sky130_fd_pr__pfet_01v8_X4L24Q_0/VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X13 a_n78_n64# a_n162_206# sky130_fd_pr__pfet_01v8_X4L24Q_0/VSUBS sky130_fd_pr__pfet_01v8_X4L24Q_0/VSUBS sky130_fd_pr__nfet_01v8 ad=0.0651 pd=0.73 as=0.0693 ps=0.75 w=0.42 l=0.15
C0 w_n260_286# a_n78_396# 3.02f
C1 a_n78_396# sky130_fd_pr__pfet_01v8_X4L24Q_0/VSUBS 2.46f
C2 w_n260_286# sky130_fd_pr__pfet_01v8_X4L24Q_0/VSUBS 6.96f
.ends

.subckt buffer_and_gate in1 clk out gnd vdd
Xbuffer_0 vdd gnd gnd gnd clk vdd m1_5444_838# vdd vdd gnd buffer
Xand_gate_0 m1_5444_838# vdd gnd in1 out and_gate
C0 in1 0 2.5f
C1 and_gate_0/a_n78_396# 0 2.34f
C2 clk 0 7.7f
C3 buffer_0/a_1436_1552# 0 8.93f
C4 vdd 0 17.7f
C5 gnd 0 7.18f
.ends

.subckt capacitor_5 m3_7768_402# buffer_and_gate_0/clk a_540_n178# a_6656_n300# w_1652_n318#
+ w_5484_n346# buffer_and_gate_0/vdd m2_n660_928# VSUBS
Xbuffer_digital_1 buffer_and_gate_0/in1 buffer_digital_1/a_116_148# buffer_and_gate_0/vdd
+ buffer_and_gate_0/vdd m2_n660_928# VSUBS VSUBS VSUBS buffer_digital
Xsky130_fd_pr__nfet_01v8_D4CMYK_0 a_6656_n300# VSUBS a_6656_n300# VSUBS VSUBS a_6656_n300#
+ VSUBS VSUBS a_6656_n300# a_6656_n300# VSUBS a_6656_n300# a_6656_n300# VSUBS a_6656_n300#
+ VSUBS VSUBS VSUBS sky130_fd_pr__nfet_01v8_D4CMYK
Xsky130_fd_pr__pfet_01v8_4ZKXAA_1 w_1652_n318# w_1652_n318# VSUBS w_1652_n318# w_1652_n318#
+ VSUBS w_1652_n318# VSUBS w_1652_n318# VSUBS VSUBS w_1652_n318# VSUBS w_1652_n318#
+ w_1652_n318# VSUBS VSUBS w_1652_n318# w_1652_n318# VSUBS w_1652_n318# VSUBS VSUBS
+ sky130_fd_pr__pfet_01v8_4ZKXAA
Xsky130_fd_pr__pfet_01v8_4ZKXAA_2 w_5484_n346# w_5484_n346# VSUBS w_5484_n346# w_5484_n346#
+ VSUBS w_5484_n346# VSUBS w_5484_n346# VSUBS VSUBS w_5484_n346# VSUBS w_5484_n346#
+ w_5484_n346# VSUBS VSUBS w_5484_n346# w_5484_n346# VSUBS w_5484_n346# VSUBS VSUBS
+ sky130_fd_pr__pfet_01v8_4ZKXAA
Xsky130_fd_pr__pfet_01v8_4ZKXAA_3 w_1652_n318# w_1652_n318# VSUBS w_1652_n318# w_1652_n318#
+ VSUBS w_1652_n318# VSUBS w_1652_n318# VSUBS VSUBS w_1652_n318# VSUBS w_1652_n318#
+ w_1652_n318# VSUBS VSUBS w_1652_n318# w_1652_n318# VSUBS w_1652_n318# VSUBS VSUBS
+ sky130_fd_pr__pfet_01v8_4ZKXAA
Xsky130_fd_pr__nfet_01v8_NJGC45_0 VSUBS a_540_n178# VSUBS a_540_n178# a_540_n178#
+ VSUBS VSUBS a_540_n178# a_540_n178# VSUBS a_540_n178# VSUBS VSUBS VSUBS VSUBS VSUBS
+ a_540_n178# VSUBS a_540_n178# a_540_n178# a_540_n178# VSUBS sky130_fd_pr__nfet_01v8_NJGC45
Xsky130_fd_pr__nfet_01v8_NJGC45_1 VSUBS w_1652_n318# VSUBS w_1652_n318# w_1652_n318#
+ VSUBS VSUBS w_1652_n318# w_1652_n318# VSUBS w_1652_n318# VSUBS VSUBS VSUBS VSUBS
+ VSUBS w_1652_n318# VSUBS w_1652_n318# w_1652_n318# w_1652_n318# VSUBS sky130_fd_pr__nfet_01v8_NJGC45
Xbuffer_and_gate_0 buffer_and_gate_0/in1 buffer_and_gate_0/clk buffer_and_gate_0/out
+ VSUBS buffer_and_gate_0/vdd buffer_and_gate
X0 buffer_and_gate_0/out m3_7768_402# sky130_fd_pr__cap_mim_m3_1 l=4.97 w=5
C0 buffer_and_gate_0/in1 m2_n660_928# 2.94f
C1 w_1652_n318# VSUBS 3.6f
C2 buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C3 buffer_and_gate_0/clk 0 7.41f
C4 buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C5 buffer_and_gate_0/vdd 0 20.2f
C6 VSUBS 0 11f
C7 a_540_n178# 0 2.32f
C8 w_1652_n318# 0 5.55f
C9 a_6656_n300# 0 2.22f
C10 buffer_and_gate_0/in1 0 2.57f
.ends

.subckt capacitors_5 m3_8778_734# capacitor_5_7/w_5484_n346# capacitor_5_7/a_6656_n300#
+ capacitor_5_7/a_540_n178# capacitor_5_5/m2_n660_928# capacitor_5_0/m2_n660_928#
+ capacitor_5_2/m2_n660_928# capacitor_5_4/m2_n660_928# capacitor_5_6/m2_n660_928#
+ capacitor_5_3/m2_n660_928# capacitor_5_7/buffer_and_gate_0/clk capacitor_5_7/w_1652_n318#
+ capacitor_5_1/m2_n660_928# capacitor_5_7/m2_n660_928# VSUBS capacitor_5_7/buffer_and_gate_0/vdd
Xcapacitor_5_5 m3_8778_734# capacitor_5_7/buffer_and_gate_0/clk capacitor_5_7/buffer_and_gate_0/vdd
+ capacitor_5_7/buffer_and_gate_0/vdd capacitor_5_7/buffer_and_gate_0/vdd capacitor_5_7/buffer_and_gate_0/vdd
+ capacitor_5_7/buffer_and_gate_0/vdd capacitor_5_5/m2_n660_928# VSUBS capacitor_5
Xcapacitor_5_6 m3_8778_734# capacitor_5_7/buffer_and_gate_0/clk capacitor_5_7/buffer_and_gate_0/vdd
+ capacitor_5_7/buffer_and_gate_0/vdd capacitor_5_7/buffer_and_gate_0/vdd capacitor_5_7/buffer_and_gate_0/vdd
+ capacitor_5_7/buffer_and_gate_0/vdd capacitor_5_6/m2_n660_928# VSUBS capacitor_5
Xcapacitor_5_7 m3_8778_734# capacitor_5_7/buffer_and_gate_0/clk capacitor_5_7/a_540_n178#
+ capacitor_5_7/a_6656_n300# capacitor_5_7/w_1652_n318# capacitor_5_7/w_5484_n346#
+ capacitor_5_7/buffer_and_gate_0/vdd capacitor_5_7/m2_n660_928# VSUBS capacitor_5
Xcapacitor_5_0 m3_8778_734# capacitor_5_7/buffer_and_gate_0/clk capacitor_5_7/buffer_and_gate_0/vdd
+ capacitor_5_7/buffer_and_gate_0/vdd capacitor_5_7/buffer_and_gate_0/vdd capacitor_5_7/buffer_and_gate_0/vdd
+ capacitor_5_7/buffer_and_gate_0/vdd capacitor_5_0/m2_n660_928# VSUBS capacitor_5
Xcapacitor_5_1 m3_8778_734# capacitor_5_7/buffer_and_gate_0/clk capacitor_5_7/buffer_and_gate_0/vdd
+ capacitor_5_7/buffer_and_gate_0/vdd capacitor_5_7/buffer_and_gate_0/vdd capacitor_5_7/buffer_and_gate_0/vdd
+ capacitor_5_7/buffer_and_gate_0/vdd capacitor_5_1/m2_n660_928# VSUBS capacitor_5
Xcapacitor_5_2 m3_8778_734# capacitor_5_7/buffer_and_gate_0/clk capacitor_5_7/buffer_and_gate_0/vdd
+ capacitor_5_7/buffer_and_gate_0/vdd capacitor_5_7/buffer_and_gate_0/vdd capacitor_5_7/buffer_and_gate_0/vdd
+ capacitor_5_7/buffer_and_gate_0/vdd capacitor_5_2/m2_n660_928# VSUBS capacitor_5
Xcapacitor_5_3 m3_8778_734# capacitor_5_7/buffer_and_gate_0/clk capacitor_5_7/buffer_and_gate_0/vdd
+ capacitor_5_7/buffer_and_gate_0/vdd capacitor_5_7/buffer_and_gate_0/vdd capacitor_5_7/buffer_and_gate_0/vdd
+ capacitor_5_7/buffer_and_gate_0/vdd capacitor_5_3/m2_n660_928# VSUBS capacitor_5
Xcapacitor_5_4 m3_8778_734# capacitor_5_7/buffer_and_gate_0/clk capacitor_5_7/buffer_and_gate_0/vdd
+ capacitor_5_7/buffer_and_gate_0/vdd capacitor_5_7/buffer_and_gate_0/vdd capacitor_5_7/buffer_and_gate_0/vdd
+ capacitor_5_7/buffer_and_gate_0/vdd capacitor_5_4/m2_n660_928# VSUBS capacitor_5
C0 capacitor_5_7/buffer_and_gate_0/clk capacitor_5_7/buffer_and_gate_0/vdd 13f
C1 VSUBS capacitor_5_7/buffer_and_gate_0/vdd 97.4f
C2 m3_8778_734# VSUBS 5.94f
C3 capacitor_5_7/buffer_and_gate_0/clk VSUBS 3.99f
C4 m3_8778_734# capacitor_5_7/buffer_and_gate_0/vdd 11.7f
C5 capacitor_5_4/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C6 capacitor_5_4/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C7 capacitor_5_4/buffer_and_gate_0/in1 0 2.57f
C8 capacitor_5_3/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C9 capacitor_5_3/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C10 capacitor_5_3/buffer_and_gate_0/in1 0 2.57f
C11 capacitor_5_2/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C12 capacitor_5_2/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C13 capacitor_5_2/buffer_and_gate_0/in1 0 2.57f
C14 capacitor_5_1/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C15 capacitor_5_1/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C16 capacitor_5_1/buffer_and_gate_0/in1 0 2.57f
C17 capacitor_5_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C18 capacitor_5_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C19 capacitor_5_0/buffer_and_gate_0/in1 0 2.57f
C20 m3_8778_734# 0 14.1f
C21 capacitor_5_7/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C22 capacitor_5_7/buffer_and_gate_0/clk 0 62.5f
C23 capacitor_5_7/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C24 capacitor_5_7/buffer_and_gate_0/vdd 0 0.18p
C25 VSUBS 0 62.2f
C26 capacitor_5_7/a_540_n178# 0 2.32f
C27 capacitor_5_7/w_1652_n318# 0 5.55f
C28 capacitor_5_7/a_6656_n300# 0 2.22f
C29 capacitor_5_7/buffer_and_gate_0/in1 0 2.57f
C30 capacitor_5_6/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C31 capacitor_5_6/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C32 capacitor_5_6/buffer_and_gate_0/in1 0 2.57f
C33 capacitor_5_5/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C34 capacitor_5_5/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C35 capacitor_5_5/buffer_and_gate_0/in1 0 2.57f
.ends

.subckt nmos_dnw3 vin out1 out2 clk clkb vs VSUBS
X0 clkb clk vin vs sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.126 ps=1.44 w=0.42 l=0.15
X1 vin clkb clk vs sky130_fd_pr__nfet_01v8 ad=0.126 pd=1.44 as=0.13 ps=1.46 w=0.42 l=0.15
X2 out2 clk vin vs sky130_fd_pr__nfet_01v8 ad=1.65 pd=7.1 as=0.945 ps=3.63 w=3 l=1
X3 vin clkb out1 vs sky130_fd_pr__nfet_01v8 ad=0.945 pd=3.63 as=1.65 ps=7.1 w=3 l=1
C0 vs VSUBS 6.64f
.ends

.subckt sky130_fd_pr__pfet_01v8_FBZ64Q a_n81_n126# a_399_n126# a_351_n223# a_n417_n223#
+ a_207_n126# a_n225_n223# a_n461_n126# a_n369_n126# a_63_157# a_303_n126# a_255_157#
+ a_n33_n223# a_15_n126# a_n177_n126# a_n129_157# a_111_n126# w_n497_n226# a_n273_n126#
+ a_159_n223# a_n321_157# VSUBS
X0 a_n273_n126# a_n321_157# a_n369_n126# w_n497_n226# sky130_fd_pr__pfet_01v8 ad=0.208 pd=1.59 as=0.208 ps=1.59 w=1.26 l=0.15
X1 a_207_n126# a_159_n223# a_111_n126# w_n497_n226# sky130_fd_pr__pfet_01v8 ad=0.208 pd=1.59 as=0.208 ps=1.59 w=1.26 l=0.15
X2 a_n177_n126# a_n225_n223# a_n273_n126# w_n497_n226# sky130_fd_pr__pfet_01v8 ad=0.208 pd=1.59 as=0.208 ps=1.59 w=1.26 l=0.15
X3 a_111_n126# a_63_157# a_15_n126# w_n497_n226# sky130_fd_pr__pfet_01v8 ad=0.208 pd=1.59 as=0.208 ps=1.59 w=1.26 l=0.15
X4 a_399_n126# a_351_n223# a_303_n126# w_n497_n226# sky130_fd_pr__pfet_01v8 ad=0.391 pd=3.14 as=0.208 ps=1.59 w=1.26 l=0.15
X5 a_n81_n126# a_n129_157# a_n177_n126# w_n497_n226# sky130_fd_pr__pfet_01v8 ad=0.208 pd=1.59 as=0.208 ps=1.59 w=1.26 l=0.15
X6 a_15_n126# a_n33_n223# a_n81_n126# w_n497_n226# sky130_fd_pr__pfet_01v8 ad=0.208 pd=1.59 as=0.208 ps=1.59 w=1.26 l=0.15
X7 a_n369_n126# a_n417_n223# a_n461_n126# w_n497_n226# sky130_fd_pr__pfet_01v8 ad=0.208 pd=1.59 as=0.391 ps=3.14 w=1.26 l=0.15
X8 a_303_n126# a_255_157# a_207_n126# w_n497_n226# sky130_fd_pr__pfet_01v8 ad=0.208 pd=1.59 as=0.208 ps=1.59 w=1.26 l=0.15
.ends

.subckt sky130_fd_pr__nfet_01v8_5ACVEW a_n129_n130# a_63_n130# a_n81_n42# a_15_n42#
+ a_n173_n42# a_n33_64# a_111_n42# VSUBS
X0 a_15_n42# a_n33_64# a_n81_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X1 a_111_n42# a_63_n130# a_15_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X2 a_n81_n42# a_n129_n130# a_n173_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
.ends

.subckt inverter_27x m1_n804_1398# m1_540_1398# m1_156_1398# m1_n36_1398# m1_732_1398#
+ m1_n1102_1398# m1_348_1398# m1_n1188_1398# m1_n996_1398# m1_n228_1398# m1_n1188_1912#
+ m1_924_1398# m1_1309_1398# a_n1158_1658# m1_n420_1398# m1_1116_1398# w_1358_2036#
+ m1_n612_1398# VSUBS
Xsky130_fd_pr__nfet_01v8_NJGLN5_1 a_n1158_1658# m1_n228_1398# a_n1158_1658# a_n1158_1658#
+ a_n1158_1658# a_n1158_1658# a_n1158_1658# m1_n1102_1398# a_n1158_1658# a_n1158_1658#
+ m1_n1102_1398# m1_n1102_1398# m1_1309_1398# m1_n420_1398# a_n1158_1658# m1_n1102_1398#
+ a_n1158_1658# a_n1158_1658# a_n1158_1658# a_n1158_1658# m1_n1102_1398# m1_540_1398#
+ m1_n1102_1398# m1_n1102_1398# a_n1158_1658# m1_n612_1398# m1_156_1398# a_n1158_1658#
+ m1_n1102_1398# a_n1158_1658# a_n1158_1658# a_n1158_1658# m1_n1102_1398# m1_732_1398#
+ a_n1158_1658# a_n1158_1658# m1_348_1398# m1_n1102_1398# m1_n804_1398# a_n1158_1658#
+ m1_924_1398# a_n1158_1658# a_n1158_1658# a_n1158_1658# a_n1158_1658# m1_n1102_1398#
+ a_n1158_1658# m1_n36_1398# m1_n1102_1398# m1_n1188_1398# m1_n996_1398# m1_n1102_1398#
+ m1_n1102_1398# m1_1116_1398# a_n1158_1658# VSUBS sky130_fd_pr__nfet_01v8_NJGLN5
Xsky130_fd_pr__pfet_01v8_VR4B8J_1 a_n1158_1658# m1_n1188_1912# m1_1309_1398# m1_1309_1398#
+ m1_n1188_1912# m1_1309_1398# a_n1158_1658# m1_1309_1398# m1_n1188_1912# a_n1158_1658#
+ a_n1158_1658# a_n1158_1658# a_n1158_1658# a_n1158_1658# a_n1158_1658# a_n1158_1658#
+ m1_n1188_1912# m1_1309_1398# m1_n1188_1912# a_n1158_1658# m1_n1188_1912# m1_n1188_1912#
+ m1_n1188_1912# a_n1158_1658# m1_1309_1398# a_n1158_1658# a_n1158_1658# a_n1158_1658#
+ a_n1158_1658# m1_1309_1398# m1_n1188_1912# a_n1158_1658# m1_n1188_1912# m1_n1188_1912#
+ a_n1158_1658# m1_n1188_1912# a_n1158_1658# w_1358_2036# m1_1309_1398# m1_1309_1398#
+ m1_1309_1398# a_n1158_1658# a_n1158_1658# a_n1158_1658# m1_1309_1398# m1_n1188_1912#
+ m1_n1188_1912# a_n1158_1658# a_n1158_1658# m1_1309_1398# a_n1158_1658# m1_1309_1398#
+ m1_1309_1398# a_n1158_1658# a_n1158_1658# a_n1158_1658# VSUBS sky130_fd_pr__pfet_01v8_VR4B8J
C0 a_n1158_1658# VSUBS 6.39f
C1 w_1358_2036# VSUBS 3.69f
.ends

.subckt sky130_fd_pr__nfet_01v8_KMMFCM a_15_n42# a_n15_n68# a_n73_n42# VSUBS
X0 a_15_n42# a_n15_n68# a_n73_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
.ends

.subckt sky130_fd_pr__pfet_01v8_29EZRJ a_n73_n126# w_n109_n188# a_15_n126# a_n15_n152#
+ VSUBS
X0 a_15_n126# a_n15_n152# a_n73_n126# w_n109_n188# sky130_fd_pr__pfet_01v8 ad=0.365 pd=3.1 as=0.365 ps=3.1 w=1.26 l=0.15
.ends

.subckt sky130_fd_pr__pfet_01v8_FL984Q a_n81_n126# a_n33_157# a_n129_n223# a_63_n223#
+ a_n173_n126# a_15_n126# a_111_n126# w_n209_n226# VSUBS
X0 a_111_n126# a_63_n223# a_15_n126# w_n209_n226# sky130_fd_pr__pfet_01v8 ad=0.391 pd=3.14 as=0.208 ps=1.59 w=1.26 l=0.15
X1 a_n81_n126# a_n129_n223# a_n173_n126# w_n209_n226# sky130_fd_pr__pfet_01v8 ad=0.208 pd=1.59 as=0.391 ps=3.14 w=1.26 l=0.15
X2 a_15_n126# a_n33_157# a_n81_n126# w_n209_n226# sky130_fd_pr__pfet_01v8 ad=0.208 pd=1.59 as=0.208 ps=1.59 w=1.26 l=0.15
.ends

.subckt sky130_fd_pr__nfet_01v8_D4CDWR a_n369_n42# a_n225_n130# a_303_n42# a_n81_n42#
+ a_399_n42# a_n33_n130# a_n273_n42# a_n461_n42# a_15_n42# a_n321_64# a_207_n42# a_159_n130#
+ a_n177_n42# a_351_n130# a_255_64# a_n417_n130# a_111_n42# a_n129_64# a_63_64# VSUBS
X0 a_303_n42# a_255_64# a_207_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X1 a_207_n42# a_159_n130# a_111_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X2 a_399_n42# a_351_n130# a_303_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X3 a_n369_n42# a_n417_n130# a_n461_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X4 a_15_n42# a_n33_n130# a_n81_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X5 a_111_n42# a_63_64# a_15_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X6 a_n273_n42# a_n321_64# a_n369_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X7 a_n81_n42# a_n129_64# a_n177_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X8 a_n177_n42# a_n225_n130# a_n273_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
.ends

.subckt clock clk_in vdd gnd clk clkb
Xsky130_fd_pr__pfet_01v8_FBZ64Q_0 vdd a_3246_118# a_2402_572# a_2402_572# a_3246_118#
+ a_2402_572# vdd a_3246_118# a_2402_572# vdd a_2402_572# a_2402_572# a_3246_118#
+ a_3246_118# a_2402_572# vdd vdd vdd a_2402_572# a_2402_572# gnd sky130_fd_pr__pfet_01v8_FBZ64Q
Xsky130_fd_pr__nfet_01v8_5ACVEW_0 a_344_n986# a_344_n986# a_2402_572# gnd gnd a_344_n986#
+ a_2402_572# gnd sky130_fd_pr__nfet_01v8_5ACVEW
Xinverter_27x_0 clk clk clk clk clk gnd clk clk clk clk vdd clk clk a_3246_118# clk
+ clk vdd clk gnd inverter_27x
Xsky130_fd_pr__nfet_01v8_KMMFCM_0 a_134_122# clk_in gnd gnd sky130_fd_pr__nfet_01v8_KMMFCM
Xsky130_fd_pr__nfet_01v8_KMMFCM_1 a_416_120# a_344_102# sky130_fd_pr__nfet_01v8_KMMFCM_2/a_15_n42#
+ gnd sky130_fd_pr__nfet_01v8_KMMFCM
Xsky130_fd_pr__nfet_01v8_KMMFCM_2 sky130_fd_pr__nfet_01v8_KMMFCM_2/a_15_n42# a_134_122#
+ gnd gnd sky130_fd_pr__nfet_01v8_KMMFCM
Xsky130_fd_pr__pfet_01v8_29EZRJ_0 vdd vdd a_134_122# clk_in gnd sky130_fd_pr__pfet_01v8_29EZRJ
Xsky130_fd_pr__pfet_01v8_FL984Q_0 a_2402_572# a_344_n986# a_344_n986# a_344_n986#
+ vdd vdd a_2402_572# vdd gnd sky130_fd_pr__pfet_01v8_FL984Q
Xsky130_fd_pr__pfet_01v8_FXZ64Q_0 vdd vdd a_1230_122# m1_998_498# gnd sky130_fd_pr__pfet_01v8_FXZ64Q
Xsky130_fd_pr__pfet_01v8_29EZRJ_1 a_416_120# vdd vdd a_344_102# gnd sky130_fd_pr__pfet_01v8_29EZRJ
Xsky130_fd_pr__pfet_01v8_FXZ64Q_1 vdd vdd a_1430_122# a_1230_122# gnd sky130_fd_pr__pfet_01v8_FXZ64Q
Xsky130_fd_pr__pfet_01v8_29EZRJ_2 vdd vdd a_416_120# a_134_122# gnd sky130_fd_pr__pfet_01v8_29EZRJ
Xsky130_fd_pr__pfet_01v8_FXZ64Q_2 vdd vdd a_344_n986# a_1430_122# gnd sky130_fd_pr__pfet_01v8_FXZ64Q
Xsky130_fd_pr__pfet_01v8_29EZRJ_3 vdd vdd m1_998_498# a_786_n2# gnd sky130_fd_pr__pfet_01v8_29EZRJ
Xsky130_fd_pr__nfet_01v8_D4CDWR_0 a_3246_118# a_2402_572# gnd gnd a_3246_118# a_2402_572#
+ gnd gnd a_3246_118# a_2402_572# a_3246_118# a_2402_572# a_3246_118# a_2402_572#
+ a_2402_572# a_2402_572# gnd a_2402_572# a_2402_572# gnd sky130_fd_pr__nfet_01v8_D4CDWR
Xsky130_fd_pr__nfet_01v8_DQBD8A_0 m1_998_498# a_786_n2# gnd gnd sky130_fd_pr__nfet_01v8_DQBD8A
Xsky130_fd_pr__nfet_01v8_DQBD8A_1 a_1230_122# m1_998_498# gnd gnd sky130_fd_pr__nfet_01v8_DQBD8A
Xsky130_fd_pr__nfet_01v8_DQBD8A_2 a_1430_122# a_1230_122# gnd gnd sky130_fd_pr__nfet_01v8_DQBD8A
Xsky130_fd_pr__nfet_01v8_DQBD8A_3 a_344_n986# a_1430_122# gnd gnd sky130_fd_pr__nfet_01v8_DQBD8A
X0 gnd a_2432_n962# clkb gnd sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X1 vdd a_2432_n962# clkb vdd sky130_fd_pr__pfet_01v8 ad=0.208 pd=1.59 as=0.208 ps=1.59 w=1.26 l=0.15
X2 vdd a_2020_n482# a_2432_n962# vdd sky130_fd_pr__pfet_01v8 ad=0.208 pd=1.59 as=0.208 ps=1.59 w=1.26 l=0.15
X3 clkb a_2432_n962# gnd gnd sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X4 vdd a_344_102# a_2020_n482# vdd sky130_fd_pr__pfet_01v8 ad=0.208 pd=1.59 as=0.208 ps=1.59 w=1.26 l=0.15
X5 gnd a_2432_n962# clkb gnd sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X6 vdd a_2432_n962# clkb vdd sky130_fd_pr__pfet_01v8 ad=0.208 pd=1.59 as=0.208 ps=1.59 w=1.26 l=0.15
X7 clkb a_2432_n962# gnd gnd sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X8 a_2020_n482# a_344_102# gnd gnd sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X9 a_786_n912# a_586_n912# vdd vdd sky130_fd_pr__pfet_01v8 ad=0.365 pd=3.1 as=0.365 ps=3.1 w=1.26 l=0.15
X10 vdd a_2432_n962# clkb vdd sky130_fd_pr__pfet_01v8 ad=0.208 pd=1.59 as=0.208 ps=1.59 w=1.26 l=0.15
X11 a_2432_n962# a_2020_n482# vdd vdd sky130_fd_pr__pfet_01v8 ad=0.208 pd=1.59 as=0.208 ps=1.59 w=1.26 l=0.15
X12 clkb a_2432_n962# vdd vdd sky130_fd_pr__pfet_01v8 ad=0.208 pd=1.59 as=0.208 ps=1.59 w=1.26 l=0.15
X13 clkb a_2432_n962# gnd gnd sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X14 gnd a_2020_n482# a_2432_n962# gnd sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X15 clkb a_2432_n962# gnd gnd sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X16 clkb a_2432_n962# vdd vdd sky130_fd_pr__pfet_01v8 ad=0.208 pd=1.59 as=0.208 ps=1.59 w=1.26 l=0.15
X17 gnd a_2432_n962# clkb gnd sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X18 gnd a_2020_n482# a_2432_n962# gnd sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X19 vdd a_2432_n962# clkb vdd sky130_fd_pr__pfet_01v8 ad=0.208 pd=1.59 as=0.208 ps=1.59 w=1.26 l=0.15
X20 a_286_n478# clk_in gnd gnd sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0.122 ps=1.42 w=0.42 l=0.15
X21 clkb a_2432_n962# vdd vdd sky130_fd_pr__pfet_01v8 ad=0.208 pd=1.59 as=0.208 ps=1.59 w=1.26 l=0.15
X22 gnd a_2432_n962# clkb gnd sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X23 a_2432_n962# a_2020_n482# vdd vdd sky130_fd_pr__pfet_01v8 ad=0.208 pd=1.59 as=0.391 ps=3.14 w=1.26 l=0.15
X24 clkb a_2432_n962# gnd gnd sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X25 a_2432_n962# a_2020_n482# gnd gnd sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X26 a_586_n2# a_416_120# gnd gnd sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X27 clkb a_2432_n962# vdd vdd sky130_fd_pr__pfet_01v8 ad=0.208 pd=1.59 as=0.208 ps=1.59 w=1.26 l=0.15
X28 gnd a_2432_n962# clkb gnd sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X29 a_2432_n962# a_2020_n482# vdd vdd sky130_fd_pr__pfet_01v8 ad=0.391 pd=3.14 as=0.208 ps=1.59 w=1.26 l=0.15
X30 a_786_n912# a_586_n912# gnd gnd sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X31 clkb a_2432_n962# vdd vdd sky130_fd_pr__pfet_01v8 ad=0.208 pd=1.59 as=0.208 ps=1.59 w=1.26 l=0.15
X32 gnd a_2432_n962# clkb gnd sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X33 vdd a_344_n986# a_286_n960# vdd sky130_fd_pr__pfet_01v8 ad=0.365 pd=3.1 as=0.183 ps=1.55 w=1.26 l=0.15
X34 a_344_102# a_1394_n918# vdd vdd sky130_fd_pr__pfet_01v8 ad=0.365 pd=3.1 as=0.365 ps=3.1 w=1.26 l=0.15
X35 a_992_n918# a_786_n912# vdd vdd sky130_fd_pr__pfet_01v8 ad=0.365 pd=3.1 as=0.365 ps=3.1 w=1.26 l=0.15
X36 a_1192_n918# a_992_n918# gnd gnd sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X37 vdd a_2432_n962# clkb vdd sky130_fd_pr__pfet_01v8 ad=0.208 pd=1.59 as=0.208 ps=1.59 w=1.26 l=0.15
X38 a_2432_n962# a_2020_n482# vdd vdd sky130_fd_pr__pfet_01v8 ad=0.208 pd=1.59 as=0.208 ps=1.59 w=1.26 l=0.15
X39 gnd a_2432_n962# clkb gnd sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X40 a_2432_n962# a_2020_n482# gnd gnd sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X41 a_1394_n918# a_1192_n918# gnd gnd sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X42 vdd a_2432_n962# clkb vdd sky130_fd_pr__pfet_01v8 ad=0.208 pd=1.59 as=0.208 ps=1.59 w=1.26 l=0.15
X43 clkb a_2432_n962# gnd gnd sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X44 clkb a_2432_n962# gnd gnd sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X45 clkb a_2432_n962# vdd vdd sky130_fd_pr__pfet_01v8 ad=0.208 pd=1.59 as=0.208 ps=1.59 w=1.26 l=0.15
X46 gnd a_2020_n482# a_2432_n962# gnd sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X47 vdd a_2432_n962# clkb vdd sky130_fd_pr__pfet_01v8 ad=0.208 pd=1.59 as=0.208 ps=1.59 w=1.26 l=0.15
X48 vdd a_2020_n482# a_2432_n962# vdd sky130_fd_pr__pfet_01v8 ad=0.208 pd=1.59 as=0.208 ps=1.59 w=1.26 l=0.15
X49 gnd a_2432_n962# clkb gnd sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X50 a_2020_n482# a_344_102# vdd vdd sky130_fd_pr__pfet_01v8 ad=0.391 pd=3.14 as=0.208 ps=1.59 w=1.26 l=0.15
X51 vdd a_2432_n962# clkb vdd sky130_fd_pr__pfet_01v8 ad=0.208 pd=1.59 as=0.208 ps=1.59 w=1.26 l=0.15
X52 clkb a_2432_n962# gnd gnd sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X53 a_586_n912# a_286_n960# vdd vdd sky130_fd_pr__pfet_01v8 ad=0.365 pd=3.1 as=0.365 ps=3.1 w=1.26 l=0.15
X54 vdd a_2020_n482# a_2432_n962# vdd sky130_fd_pr__pfet_01v8 ad=0.208 pd=1.59 as=0.208 ps=1.59 w=1.26 l=0.15
X55 a_586_n2# a_416_120# vdd vdd sky130_fd_pr__pfet_01v8 ad=0.365 pd=3.1 as=0.365 ps=3.1 w=1.26 l=0.15
X56 clkb a_2432_n962# vdd vdd sky130_fd_pr__pfet_01v8 ad=0.208 pd=1.59 as=0.391 ps=3.14 w=1.26 l=0.15
X57 clkb a_2432_n962# vdd vdd sky130_fd_pr__pfet_01v8 ad=0.208 pd=1.59 as=0.208 ps=1.59 w=1.26 l=0.15
X58 vdd a_2432_n962# clkb vdd sky130_fd_pr__pfet_01v8 ad=0.208 pd=1.59 as=0.208 ps=1.59 w=1.26 l=0.15
X59 clkb a_2432_n962# gnd gnd sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X60 gnd a_2432_n962# clkb gnd sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X61 gnd a_2020_n482# a_2432_n962# gnd sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X62 clkb a_2432_n962# vdd vdd sky130_fd_pr__pfet_01v8 ad=0.208 pd=1.59 as=0.208 ps=1.59 w=1.26 l=0.15
X63 gnd a_2432_n962# clkb gnd sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X64 clkb a_2432_n962# gnd gnd sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X65 clkb a_2432_n962# vdd vdd sky130_fd_pr__pfet_01v8 ad=0.208 pd=1.59 as=0.208 ps=1.59 w=1.26 l=0.15
X66 a_2020_n482# a_344_102# gnd gnd sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X67 vdd a_2432_n962# clkb vdd sky130_fd_pr__pfet_01v8 ad=0.208 pd=1.59 as=0.208 ps=1.59 w=1.26 l=0.15
X68 gnd a_2432_n962# clkb gnd sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X69 a_2432_n962# a_2020_n482# gnd gnd sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X70 gnd a_2432_n962# clkb gnd sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X71 a_786_n2# a_586_n2# gnd gnd sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X72 clkb a_2432_n962# gnd gnd sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X73 a_286_n960# clk_in vdd vdd sky130_fd_pr__pfet_01v8 ad=0.183 pd=1.55 as=0.365 ps=3.1 w=1.26 l=0.15
X74 clkb a_2432_n962# vdd vdd sky130_fd_pr__pfet_01v8 ad=0.208 pd=1.59 as=0.208 ps=1.59 w=1.26 l=0.15
X75 a_286_n960# a_344_n986# a_286_n478# gnd sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0609 ps=0.71 w=0.42 l=0.15
X76 a_2432_n962# a_2020_n482# vdd vdd sky130_fd_pr__pfet_01v8 ad=0.208 pd=1.59 as=0.208 ps=1.59 w=1.26 l=0.15
X77 a_586_n912# a_286_n960# gnd gnd sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X78 a_1394_n918# a_1192_n918# vdd vdd sky130_fd_pr__pfet_01v8 ad=0.365 pd=3.1 as=0.365 ps=3.1 w=1.26 l=0.15
X79 a_1192_n918# a_992_n918# vdd vdd sky130_fd_pr__pfet_01v8 ad=0.365 pd=3.1 as=0.365 ps=3.1 w=1.26 l=0.15
X80 gnd a_2432_n962# clkb gnd sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X81 a_2432_n962# a_2020_n482# gnd gnd sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X82 vdd a_2432_n962# clkb vdd sky130_fd_pr__pfet_01v8 ad=0.208 pd=1.59 as=0.208 ps=1.59 w=1.26 l=0.15
X83 clkb a_2432_n962# vdd vdd sky130_fd_pr__pfet_01v8 ad=0.208 pd=1.59 as=0.208 ps=1.59 w=1.26 l=0.15
X84 vdd a_2020_n482# a_2432_n962# vdd sky130_fd_pr__pfet_01v8 ad=0.208 pd=1.59 as=0.208 ps=1.59 w=1.26 l=0.15
X85 vdd a_2432_n962# clkb vdd sky130_fd_pr__pfet_01v8 ad=0.208 pd=1.59 as=0.208 ps=1.59 w=1.26 l=0.15
X86 a_2432_n962# a_2020_n482# gnd gnd sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X87 a_344_102# a_1394_n918# gnd gnd sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X88 a_2020_n482# a_344_102# vdd vdd sky130_fd_pr__pfet_01v8 ad=0.208 pd=1.59 as=0.391 ps=3.14 w=1.26 l=0.15
X89 clkb a_2432_n962# gnd gnd sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X90 gnd a_344_102# a_2020_n482# gnd sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X91 a_992_n918# a_786_n912# gnd gnd sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X92 gnd a_2432_n962# clkb gnd sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X93 clkb a_2432_n962# vdd vdd sky130_fd_pr__pfet_01v8 ad=0.391 pd=3.14 as=0.208 ps=1.59 w=1.26 l=0.15
X94 vdd a_2432_n962# clkb vdd sky130_fd_pr__pfet_01v8 ad=0.208 pd=1.59 as=0.208 ps=1.59 w=1.26 l=0.15
X95 clkb a_2432_n962# gnd gnd sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X96 a_786_n2# a_586_n2# vdd vdd sky130_fd_pr__pfet_01v8 ad=0.365 pd=3.1 as=0.365 ps=3.1 w=1.26 l=0.15
X97 clkb a_2432_n962# vdd vdd sky130_fd_pr__pfet_01v8 ad=0.208 pd=1.59 as=0.208 ps=1.59 w=1.26 l=0.15
C0 vdd clkb 7.31f
C1 vdd a_2432_n962# 7.04f
C2 clkb a_2432_n962# 2.67f
C3 a_2020_n482# vdd 2.66f
C4 clkb gnd 5.1f
C5 a_2432_n962# gnd 8.71f
C6 a_2020_n482# gnd 2.57f
C7 vdd gnd 26.1f
C8 a_344_102# gnd 2.81f
C9 a_2402_572# gnd 2.31f
C10 a_344_n986# gnd 2.43f
C11 a_3246_118# gnd 6.79f
.ends

.subckt sky130_fd_pr__pfet_01v8_4RPJ49 a_2031_73# a_1887_n42# a_3615_n42# a_3183_73#
+ a_n3729_73# a_n2529_n42# a_1503_n42# a_63_n42# a_n753_n139# a_n3393_n42# a_n369_n139#
+ a_n1425_73# a_n1281_n42# a_n2961_73# a_687_73# a_n2577_73# a_n417_n42# a_2367_n42#
+ a_n1761_n42# a_n3009_n42# a_n2673_n139# a_2847_n42# a_n2289_n139# a_n3633_n139#
+ a_2607_73# a_n3249_n139# a_n1713_n139# a_3759_73# a_n1329_n139# a_255_n42# a_1455_73#
+ a_n2241_n42# a_2991_73# a_3471_n139# a_735_n42# a_1551_n139# a_3087_n139# a_1599_n42#
+ a_3327_n42# a_1167_n139# a_n2721_n42# a_n81_73# a_2511_n139# a_1215_n42# a_n273_73#
+ a_2127_n139# a_n993_n42# a_3807_n42# a_15_n139# a_303_73# a_n3585_n42# a_n129_n42#
+ a_2079_n42# a_n561_n139# a_n3345_73# a_n3201_n42# a_n1473_n42# a_n177_n139# a_n1041_73#
+ a_n609_n42# a_2559_n42# a_n2193_73# a_n1953_n42# a_n849_73# w_n3905_n142# a_n2481_n139#
+ a_n2097_n139# a_n3441_n139# a_1791_n42# a_n1521_n139# a_n3057_n139# a_2223_73# a_447_n42#
+ a_3039_n42# a_n1137_n139# a_3375_73# a_n2433_n42# a_927_n42# a_1071_73# a_n1617_73#
+ a_n2913_n42# a_3519_n42# a_975_n139# a_879_73# a_n2769_73# a_n321_n42# a_1407_n42#
+ a_n3297_n42# a_2271_n42# a_n1185_n42# a_n801_n42# a_n3777_n42# a_2751_n42# a_n1665_n42#
+ a_1647_73# a_2799_73# a_3231_n42# a_159_n42# a_n2145_n42# a_n465_73# a_1983_n42#
+ a_3711_n42# a_639_n42# a_n2625_n42# a_1119_n42# a_n3537_73# a_n897_n42# a_n513_n42#
+ a_n1233_73# a_n3489_n42# a_2463_n42# a_783_n139# a_495_73# a_399_n139# a_n2385_73#
+ a_2895_n139# a_n3105_n42# a_n1377_n42# a_2943_n42# a_1935_n139# a_n1857_n42# a_351_n42#
+ a_2415_73# a_n33_n42# a_3567_73# a_831_n42# a_1695_n42# a_3423_n42# a_1263_73# a_n945_n139#
+ a_n2337_n42# a_1311_n42# a_n1809_73# a_n2817_n42# a_n3681_n42# a_n225_n42# a_2175_n42#
+ a_n2865_n139# a_n1089_n42# a_n3825_n139# a_111_73# a_n2001_73# a_n3869_n42# a_n705_n42#
+ a_2655_n42# a_n1905_n139# a_n3153_73# a_591_n139# a_1839_73# a_n1569_n42# a_3663_n139#
+ a_1743_n139# a_3279_n139# a_543_n42# a_207_n139# a_n657_73# a_1359_n139# a_2703_n139#
+ a_3135_n42# VSUBS a_2319_n139# a_n2049_n42# a_1023_n42#
X0 a_n2241_n42# a_n2289_n139# a_n2337_n42# w_n3905_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X1 a_n2913_n42# a_n2961_73# a_n3009_n42# w_n3905_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X2 a_n2721_n42# a_n2769_73# a_n2817_n42# w_n3905_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X3 a_n2625_n42# a_n2673_n139# a_n2721_n42# w_n3905_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X4 a_n2433_n42# a_n2481_n139# a_n2529_n42# w_n3905_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X5 a_n2337_n42# a_n2385_73# a_n2433_n42# w_n3905_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X6 a_n2145_n42# a_n2193_73# a_n2241_n42# w_n3905_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X7 a_n2049_n42# a_n2097_n139# a_n2145_n42# w_n3905_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X8 a_n2817_n42# a_n2865_n139# a_n2913_n42# w_n3905_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X9 a_n2529_n42# a_n2577_73# a_n2625_n42# w_n3905_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X10 a_2079_n42# a_2031_73# a_1983_n42# w_n3905_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X11 a_2175_n42# a_2127_n139# a_2079_n42# w_n3905_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X12 a_2271_n42# a_2223_73# a_2175_n42# w_n3905_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X13 a_2367_n42# a_2319_n139# a_2271_n42# w_n3905_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X14 a_2463_n42# a_2415_73# a_2367_n42# w_n3905_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X15 a_2655_n42# a_2607_73# a_2559_n42# w_n3905_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X16 a_2751_n42# a_2703_n139# a_2655_n42# w_n3905_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X17 a_2943_n42# a_2895_n139# a_2847_n42# w_n3905_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X18 a_2559_n42# a_2511_n139# a_2463_n42# w_n3905_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X19 a_2847_n42# a_2799_73# a_2751_n42# w_n3905_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X20 a_927_n42# a_879_73# a_831_n42# w_n3905_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X21 a_1023_n42# a_975_n139# a_927_n42# w_n3905_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X22 a_n1953_n42# a_n2001_73# a_n2049_n42# w_n3905_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X23 a_n1761_n42# a_n1809_73# a_n1857_n42# w_n3905_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X24 a_n1665_n42# a_n1713_n139# a_n1761_n42# w_n3905_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X25 a_n1857_n42# a_n1905_n139# a_n1953_n42# w_n3905_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X26 a_n1569_n42# a_n1617_73# a_n1665_n42# w_n3905_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X27 a_1119_n42# a_1071_73# a_1023_n42# w_n3905_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X28 a_1215_n42# a_1167_n139# a_1119_n42# w_n3905_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X29 a_1311_n42# a_1263_73# a_1215_n42# w_n3905_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X30 a_1407_n42# a_1359_n139# a_1311_n42# w_n3905_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X31 a_1503_n42# a_1455_73# a_1407_n42# w_n3905_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X32 a_1695_n42# a_1647_73# a_1599_n42# w_n3905_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X33 a_1791_n42# a_1743_n139# a_1695_n42# w_n3905_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X34 a_1599_n42# a_1551_n139# a_1503_n42# w_n3905_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X35 a_1887_n42# a_1839_73# a_1791_n42# w_n3905_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X36 a_1983_n42# a_1935_n139# a_1887_n42# w_n3905_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X37 a_n33_n42# a_n81_73# a_n129_n42# w_n3905_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X38 a_351_n42# a_303_73# a_255_n42# w_n3905_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X39 a_159_n42# a_111_73# a_63_n42# w_n3905_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X40 a_255_n42# a_207_n139# a_159_n42# w_n3905_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X41 a_447_n42# a_399_n139# a_351_n42# w_n3905_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X42 a_543_n42# a_495_73# a_447_n42# w_n3905_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X43 a_639_n42# a_591_n139# a_543_n42# w_n3905_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X44 a_735_n42# a_687_73# a_639_n42# w_n3905_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X45 a_831_n42# a_783_n139# a_735_n42# w_n3905_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X46 a_n1473_n42# a_n1521_n139# a_n1569_n42# w_n3905_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X47 a_n1377_n42# a_n1425_73# a_n1473_n42# w_n3905_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X48 a_n1281_n42# a_n1329_n139# a_n1377_n42# w_n3905_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X49 a_n1185_n42# a_n1233_73# a_n1281_n42# w_n3905_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X50 a_n1089_n42# a_n1137_n139# a_n1185_n42# w_n3905_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X51 a_n993_n42# a_n1041_73# a_n1089_n42# w_n3905_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X52 a_n801_n42# a_n849_73# a_n897_n42# w_n3905_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X53 a_n513_n42# a_n561_n139# a_n609_n42# w_n3905_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X54 a_n321_n42# a_n369_n139# a_n417_n42# w_n3905_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X55 a_n225_n42# a_n273_73# a_n321_n42# w_n3905_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X56 a_n897_n42# a_n945_n139# a_n993_n42# w_n3905_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X57 a_n705_n42# a_n753_n139# a_n801_n42# w_n3905_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X58 a_n609_n42# a_n657_73# a_n705_n42# w_n3905_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X59 a_n417_n42# a_n465_73# a_n513_n42# w_n3905_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X60 a_n129_n42# a_n177_n139# a_n225_n42# w_n3905_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X61 a_3327_n42# a_3279_n139# a_3231_n42# w_n3905_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X62 a_3423_n42# a_3375_73# a_3327_n42# w_n3905_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X63 a_3615_n42# a_3567_73# a_3519_n42# w_n3905_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X64 a_3711_n42# a_3663_n139# a_3615_n42# w_n3905_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X65 a_3519_n42# a_3471_n139# a_3423_n42# w_n3905_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X66 a_3807_n42# a_3759_73# a_3711_n42# w_n3905_n142# sky130_fd_pr__pfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X67 a_n3201_n42# a_n3249_n139# a_n3297_n42# w_n3905_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X68 a_63_n42# a_15_n139# a_n33_n42# w_n3905_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X69 a_n3681_n42# a_n3729_73# a_n3777_n42# w_n3905_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X70 a_n3585_n42# a_n3633_n139# a_n3681_n42# w_n3905_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X71 a_n3393_n42# a_n3441_n139# a_n3489_n42# w_n3905_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X72 a_n3297_n42# a_n3345_73# a_n3393_n42# w_n3905_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X73 a_n3105_n42# a_n3153_73# a_n3201_n42# w_n3905_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X74 a_n3009_n42# a_n3057_n139# a_n3105_n42# w_n3905_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X75 a_3231_n42# a_3183_73# a_3135_n42# w_n3905_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X76 a_n3777_n42# a_n3825_n139# a_n3869_n42# w_n3905_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X77 a_n3489_n42# a_n3537_73# a_n3585_n42# w_n3905_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X78 a_3039_n42# a_2991_73# a_2943_n42# w_n3905_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X79 a_3135_n42# a_3087_n139# a_3039_n42# w_n3905_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
C0 w_n3905_n142# VSUBS 6.63f
.ends

.subckt sky130_fd_pr__nfet_01v8_NJGC8F a_15_n130# a_1887_n42# a_3615_n42# a_1647_64#
+ a_n561_n130# a_n2529_n42# a_1503_n42# a_2799_64# a_63_n42# a_n177_n130# a_n3393_n42#
+ a_n1281_n42# a_n465_64# a_n417_n42# a_2367_n42# a_n1761_n42# a_n2481_n130# a_n3009_n42#
+ a_n2097_n130# a_n3441_n130# a_2847_n42# a_n1521_n130# a_n3057_n130# a_n3537_64#
+ a_n1137_n130# a_255_n42# a_n1233_64# a_495_64# a_n2241_n42# a_n2385_64# a_975_n130#
+ a_735_n42# a_1599_n42# a_3327_n42# a_n2721_n42# a_1215_n42# a_2415_64# a_n993_n42#
+ a_3807_n42# a_3567_64# a_n3585_n42# a_n129_n42# a_2079_n42# a_1263_64# a_n3201_n42#
+ a_n1473_n42# a_n1809_64# a_n609_n42# a_2559_n42# a_n1953_n42# a_111_64# a_n2001_64#
+ a_1791_n42# a_447_n42# a_n3153_64# a_3039_n42# a_n2433_n42# a_1839_64# a_927_n42#
+ a_n2913_n42# a_3519_n42# a_783_n130# a_399_n130# a_2895_n130# a_n321_n42# a_1407_n42#
+ a_n3297_n42# a_2271_n42# a_n657_64# a_n1185_n42# a_1935_n130# a_n801_n42# a_2031_64#
+ a_n3777_n42# a_2751_n42# a_3183_64# a_n1665_n42# a_n3729_64# a_n1425_64# a_687_64#
+ a_n2961_64# a_n945_n130# a_n2577_64# a_3231_n42# a_159_n42# a_n2145_n42# a_1983_n42#
+ a_3711_n42# a_2607_64# a_639_n42# a_n2625_n42# a_3759_64# a_n2865_n130# a_1119_n42#
+ a_n3825_n130# a_1455_64# a_n1905_n130# a_2991_64# a_n897_n42# a_591_n130# a_n513_n42#
+ a_n3489_n42# a_2463_n42# a_n3105_n42# a_n1377_n42# a_n81_64# a_n273_64# a_3663_n130#
+ a_3279_n130# a_2943_n42# a_1743_n130# a_207_n130# a_2703_n130# a_1359_n130# a_n1857_n42#
+ a_2319_n130# a_351_n42# a_303_64# a_n3345_64# a_n33_n42# a_831_n42# a_n1041_64#
+ a_1695_n42# a_3423_n42# a_n753_n130# a_n369_n130# a_n2193_64# a_n2337_n42# a_1311_n42#
+ a_n849_64# a_n2817_n42# a_n3681_n42# a_n225_n42# a_2223_64# a_n2673_n130# a_2175_n42#
+ a_3375_64# a_n2289_n130# a_n3633_n130# a_n1089_n42# a_n3249_n130# a_n1713_n130#
+ a_n3869_n42# a_n705_n42# a_2655_n42# a_1071_64# a_n1329_n130# a_n1617_64# a_n1569_n42#
+ a_879_64# a_n2769_64# a_3471_n130# a_3087_n130# a_1551_n130# a_2511_n130# a_543_n42#
+ a_1167_n130# a_3135_n42# a_2127_n130# VSUBS a_n2049_n42# a_1023_n42#
X0 a_n3201_n42# a_n3249_n130# a_n3297_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X1 a_63_n42# a_15_n130# a_n33_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X2 a_n3681_n42# a_n3729_64# a_n3777_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X3 a_n3585_n42# a_n3633_n130# a_n3681_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X4 a_n3393_n42# a_n3441_n130# a_n3489_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X5 a_n3297_n42# a_n3345_64# a_n3393_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X6 a_n3105_n42# a_n3153_64# a_n3201_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X7 a_n3009_n42# a_n3057_n130# a_n3105_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X8 a_n3777_n42# a_n3825_n130# a_n3869_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X9 a_n3489_n42# a_n3537_64# a_n3585_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X10 a_3135_n42# a_3087_n130# a_3039_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X11 a_3231_n42# a_3183_64# a_3135_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X12 a_3039_n42# a_2991_64# a_2943_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X13 a_n2241_n42# a_n2289_n130# a_n2337_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X14 a_n2913_n42# a_n2961_64# a_n3009_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X15 a_n2721_n42# a_n2769_64# a_n2817_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X16 a_n2625_n42# a_n2673_n130# a_n2721_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X17 a_n2433_n42# a_n2481_n130# a_n2529_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X18 a_n2337_n42# a_n2385_64# a_n2433_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X19 a_n2145_n42# a_n2193_64# a_n2241_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X20 a_n2049_n42# a_n2097_n130# a_n2145_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X21 a_n2817_n42# a_n2865_n130# a_n2913_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X22 a_n2529_n42# a_n2577_64# a_n2625_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X23 a_2175_n42# a_2127_n130# a_2079_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X24 a_2271_n42# a_2223_64# a_2175_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X25 a_2463_n42# a_2415_64# a_2367_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X26 a_2751_n42# a_2703_n130# a_2655_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X27 a_2079_n42# a_2031_64# a_1983_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X28 a_2367_n42# a_2319_n130# a_2271_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X29 a_2559_n42# a_2511_n130# a_2463_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X30 a_2655_n42# a_2607_64# a_2559_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X31 a_2847_n42# a_2799_64# a_2751_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X32 a_2943_n42# a_2895_n130# a_2847_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X33 a_927_n42# a_879_64# a_831_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X34 a_1023_n42# a_975_n130# a_927_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X35 a_n1953_n42# a_n2001_64# a_n2049_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X36 a_n1761_n42# a_n1809_64# a_n1857_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X37 a_n1665_n42# a_n1713_n130# a_n1761_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X38 a_n1857_n42# a_n1905_n130# a_n1953_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X39 a_n1569_n42# a_n1617_64# a_n1665_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X40 a_1215_n42# a_1167_n130# a_1119_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X41 a_1311_n42# a_1263_64# a_1215_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X42 a_1503_n42# a_1455_64# a_1407_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X43 a_1791_n42# a_1743_n130# a_1695_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X44 a_1119_n42# a_1071_64# a_1023_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X45 a_1407_n42# a_1359_n130# a_1311_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X46 a_1599_n42# a_1551_n130# a_1503_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X47 a_1695_n42# a_1647_64# a_1599_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X48 a_1887_n42# a_1839_64# a_1791_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X49 a_1983_n42# a_1935_n130# a_1887_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X50 a_n33_n42# a_n81_64# a_n129_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X51 a_351_n42# a_303_64# a_255_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X52 a_159_n42# a_111_64# a_63_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X53 a_255_n42# a_207_n130# a_159_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X54 a_447_n42# a_399_n130# a_351_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X55 a_543_n42# a_495_64# a_447_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X56 a_735_n42# a_687_64# a_639_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X57 a_831_n42# a_783_n130# a_735_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X58 a_639_n42# a_591_n130# a_543_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X59 a_n1473_n42# a_n1521_n130# a_n1569_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X60 a_n1281_n42# a_n1329_n130# a_n1377_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X61 a_n1185_n42# a_n1233_64# a_n1281_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X62 a_n993_n42# a_n1041_64# a_n1089_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X63 a_n1377_n42# a_n1425_64# a_n1473_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X64 a_n1089_n42# a_n1137_n130# a_n1185_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X65 a_n321_n42# a_n369_n130# a_n417_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X66 a_n801_n42# a_n849_64# a_n897_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X67 a_n705_n42# a_n753_n130# a_n801_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X68 a_n609_n42# a_n657_64# a_n705_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X69 a_n513_n42# a_n561_n130# a_n609_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X70 a_n417_n42# a_n465_64# a_n513_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X71 a_n225_n42# a_n273_64# a_n321_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X72 a_n129_n42# a_n177_n130# a_n225_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X73 a_n897_n42# a_n945_n130# a_n993_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X74 a_3327_n42# a_3279_n130# a_3231_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X75 a_3423_n42# a_3375_64# a_3327_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X76 a_3615_n42# a_3567_64# a_3519_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X77 a_3711_n42# a_3663_n130# a_3615_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X78 a_3519_n42# a_3471_n130# a_3423_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X79 a_3807_n42# a_3759_64# a_3711_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
.ends

.subckt nmos_diode2 a_350_n764# a_970_n762# a_410_n892# dw_118_n1078# VSUBS
X0 a_410_n892# a_410_n892# a_350_n764# dw_118_n1078# sky130_fd_pr__nfet_01v8 ad=0.873 pd=6.6 as=0.903 ps=6.62 w=3.01 l=1
X1 a_350_n764# a_970_n762# a_970_n762# dw_118_n1078# sky130_fd_pr__nfet_01v8 ad=0.993 pd=6.68 as=0.873 ps=6.6 w=3.01 l=1
C0 dw_118_n1078# VSUBS 8.16f
.ends

.subckt charge_pump m1_12174_n760# nmos_dnw3_0/vin m2_10426_9616# clock_0/clk_in m2_10400_5448#
+ m2_10388_7530# m2_10266_15868# m2_10336_11702# m2_10436_1276# m2_10362_3360# m2_10308_13784#
+ clock_0/vdd nmos_dnw3_0/vs clock_0/gnd
Xsky130_fd_pr__cap_mim_m3_1_MH6KF8_4 nmos_dnw3_0/clk clock_0/clk clock_0/gnd sky130_fd_pr__cap_mim_m3_1_MH6KF8
Xsky130_fd_pr__cap_mim_m3_1_MH6KF8_5 nmos_dnw3_0/clkb clock_0/clkb clock_0/gnd sky130_fd_pr__cap_mim_m3_1_MH6KF8
Xcapacitors_5_1 nmos_dnw3_0/out2 clock_0/vdd clock_0/vdd clock_0/vdd m2_10400_5448#
+ m2_10266_15868# m2_10336_11702# m2_10388_7530# m2_10362_3360# m2_10426_9616# clock_0/clkb
+ clock_0/vdd m2_10308_13784# m2_10436_1276# clock_0/gnd clock_0/vdd capacitors_5
Xcapacitors_5_0 nmos_dnw3_0/out1 clock_0/vdd clock_0/vdd clock_0/vdd m2_10400_5448#
+ m2_10266_15868# m2_10336_11702# m2_10388_7530# m2_10362_3360# m2_10426_9616# clock_0/clk
+ clock_0/vdd m2_10308_13784# m2_10436_1276# clock_0/gnd clock_0/vdd capacitors_5
Xnmos_dnw3_0 nmos_dnw3_0/vin nmos_dnw3_0/out1 nmos_dnw3_0/out2 nmos_dnw3_0/clk nmos_dnw3_0/clkb
+ nmos_dnw3_0/vs clock_0/gnd nmos_dnw3
Xclock_0 clock_0/clk_in clock_0/vdd clock_0/gnd clock_0/clk clock_0/clkb clock
Xsky130_fd_pr__pfet_01v8_4RPJ49_0 clock_0/gnd clock_0/vdd clock_0/vdd clock_0/gnd
+ clock_0/gnd clock_0/vdd clock_0/vdd clock_0/vdd clock_0/gnd clock_0/vdd clock_0/gnd
+ clock_0/gnd clock_0/vdd clock_0/gnd clock_0/gnd clock_0/gnd clock_0/vdd clock_0/vdd
+ clock_0/vdd clock_0/vdd clock_0/gnd clock_0/vdd clock_0/gnd clock_0/gnd clock_0/gnd
+ clock_0/gnd clock_0/gnd clock_0/gnd clock_0/gnd clock_0/vdd clock_0/gnd clock_0/vdd
+ clock_0/gnd clock_0/gnd clock_0/vdd clock_0/gnd clock_0/gnd clock_0/vdd clock_0/vdd
+ clock_0/gnd clock_0/vdd clock_0/gnd clock_0/gnd clock_0/vdd clock_0/gnd clock_0/gnd
+ clock_0/vdd clock_0/vdd clock_0/gnd clock_0/gnd clock_0/vdd clock_0/vdd clock_0/vdd
+ clock_0/gnd clock_0/gnd clock_0/vdd clock_0/vdd clock_0/gnd clock_0/gnd clock_0/vdd
+ clock_0/vdd clock_0/gnd clock_0/vdd clock_0/gnd clock_0/vdd clock_0/gnd clock_0/gnd
+ clock_0/gnd clock_0/vdd clock_0/gnd clock_0/gnd clock_0/gnd clock_0/vdd clock_0/vdd
+ clock_0/gnd clock_0/gnd clock_0/vdd clock_0/vdd clock_0/gnd clock_0/gnd clock_0/vdd
+ clock_0/vdd clock_0/gnd clock_0/gnd clock_0/gnd clock_0/vdd clock_0/vdd clock_0/vdd
+ clock_0/vdd clock_0/vdd clock_0/vdd clock_0/vdd clock_0/vdd clock_0/vdd clock_0/gnd
+ clock_0/gnd clock_0/vdd clock_0/vdd clock_0/vdd clock_0/gnd clock_0/vdd clock_0/vdd
+ clock_0/vdd clock_0/vdd clock_0/vdd clock_0/gnd clock_0/vdd clock_0/vdd clock_0/gnd
+ clock_0/vdd clock_0/vdd clock_0/gnd clock_0/gnd clock_0/gnd clock_0/gnd clock_0/gnd
+ clock_0/vdd clock_0/vdd clock_0/vdd clock_0/gnd clock_0/vdd clock_0/vdd clock_0/gnd
+ clock_0/vdd clock_0/gnd clock_0/vdd clock_0/vdd clock_0/vdd clock_0/gnd clock_0/gnd
+ clock_0/vdd clock_0/vdd clock_0/gnd clock_0/vdd clock_0/vdd clock_0/vdd clock_0/vdd
+ clock_0/gnd clock_0/vdd clock_0/gnd clock_0/gnd clock_0/gnd clock_0/vdd clock_0/vdd
+ clock_0/vdd clock_0/gnd clock_0/gnd clock_0/gnd clock_0/gnd clock_0/vdd clock_0/gnd
+ clock_0/gnd clock_0/gnd clock_0/vdd clock_0/gnd clock_0/gnd clock_0/gnd clock_0/gnd
+ clock_0/vdd clock_0/gnd clock_0/gnd clock_0/vdd clock_0/vdd sky130_fd_pr__pfet_01v8_4RPJ49
Xsky130_fd_pr__pfet_01v8_4RPJ49_1 clock_0/gnd clock_0/vdd clock_0/vdd clock_0/gnd
+ clock_0/gnd clock_0/vdd clock_0/vdd clock_0/vdd clock_0/gnd clock_0/vdd clock_0/gnd
+ clock_0/gnd clock_0/vdd clock_0/gnd clock_0/gnd clock_0/gnd clock_0/vdd clock_0/vdd
+ clock_0/vdd clock_0/vdd clock_0/gnd clock_0/vdd clock_0/gnd clock_0/gnd clock_0/gnd
+ clock_0/gnd clock_0/gnd clock_0/gnd clock_0/gnd clock_0/vdd clock_0/gnd clock_0/vdd
+ clock_0/gnd clock_0/gnd clock_0/vdd clock_0/gnd clock_0/gnd clock_0/vdd clock_0/vdd
+ clock_0/gnd clock_0/vdd clock_0/gnd clock_0/gnd clock_0/vdd clock_0/gnd clock_0/gnd
+ clock_0/vdd clock_0/vdd clock_0/gnd clock_0/gnd clock_0/vdd clock_0/vdd clock_0/vdd
+ clock_0/gnd clock_0/gnd clock_0/vdd clock_0/vdd clock_0/gnd clock_0/gnd clock_0/vdd
+ clock_0/vdd clock_0/gnd clock_0/vdd clock_0/gnd clock_0/vdd clock_0/gnd clock_0/gnd
+ clock_0/gnd clock_0/vdd clock_0/gnd clock_0/gnd clock_0/gnd clock_0/vdd clock_0/vdd
+ clock_0/gnd clock_0/gnd clock_0/vdd clock_0/vdd clock_0/gnd clock_0/gnd clock_0/vdd
+ clock_0/vdd clock_0/gnd clock_0/gnd clock_0/gnd clock_0/vdd clock_0/vdd clock_0/vdd
+ clock_0/vdd clock_0/vdd clock_0/vdd clock_0/vdd clock_0/vdd clock_0/vdd clock_0/gnd
+ clock_0/gnd clock_0/vdd clock_0/vdd clock_0/vdd clock_0/gnd clock_0/vdd clock_0/vdd
+ clock_0/vdd clock_0/vdd clock_0/vdd clock_0/gnd clock_0/vdd clock_0/vdd clock_0/gnd
+ clock_0/vdd clock_0/vdd clock_0/gnd clock_0/gnd clock_0/gnd clock_0/gnd clock_0/gnd
+ clock_0/vdd clock_0/vdd clock_0/vdd clock_0/gnd clock_0/vdd clock_0/vdd clock_0/gnd
+ clock_0/vdd clock_0/gnd clock_0/vdd clock_0/vdd clock_0/vdd clock_0/gnd clock_0/gnd
+ clock_0/vdd clock_0/vdd clock_0/gnd clock_0/vdd clock_0/vdd clock_0/vdd clock_0/vdd
+ clock_0/gnd clock_0/vdd clock_0/gnd clock_0/gnd clock_0/gnd clock_0/vdd clock_0/vdd
+ clock_0/vdd clock_0/gnd clock_0/gnd clock_0/gnd clock_0/gnd clock_0/vdd clock_0/gnd
+ clock_0/gnd clock_0/gnd clock_0/vdd clock_0/gnd clock_0/gnd clock_0/gnd clock_0/gnd
+ clock_0/vdd clock_0/gnd clock_0/gnd clock_0/vdd clock_0/vdd sky130_fd_pr__pfet_01v8_4RPJ49
Xsky130_fd_pr__nfet_01v8_NJGC8F_0 clock_0/vdd clock_0/gnd clock_0/gnd clock_0/vdd
+ clock_0/vdd clock_0/gnd clock_0/gnd clock_0/vdd clock_0/gnd clock_0/vdd clock_0/gnd
+ clock_0/gnd clock_0/vdd clock_0/gnd clock_0/gnd clock_0/gnd clock_0/vdd clock_0/gnd
+ clock_0/vdd clock_0/vdd clock_0/gnd clock_0/vdd clock_0/vdd clock_0/vdd clock_0/vdd
+ clock_0/gnd clock_0/vdd clock_0/vdd clock_0/gnd clock_0/vdd clock_0/vdd clock_0/gnd
+ clock_0/gnd clock_0/gnd clock_0/gnd clock_0/gnd clock_0/vdd clock_0/gnd clock_0/gnd
+ clock_0/vdd clock_0/gnd clock_0/gnd clock_0/gnd clock_0/vdd clock_0/gnd clock_0/gnd
+ clock_0/vdd clock_0/gnd clock_0/gnd clock_0/gnd clock_0/vdd clock_0/vdd clock_0/gnd
+ clock_0/gnd clock_0/vdd clock_0/gnd clock_0/gnd clock_0/vdd clock_0/gnd clock_0/gnd
+ clock_0/gnd clock_0/vdd clock_0/vdd clock_0/vdd clock_0/gnd clock_0/gnd clock_0/gnd
+ clock_0/gnd clock_0/vdd clock_0/gnd clock_0/vdd clock_0/gnd clock_0/vdd clock_0/gnd
+ clock_0/gnd clock_0/vdd clock_0/gnd clock_0/vdd clock_0/vdd clock_0/vdd clock_0/vdd
+ clock_0/vdd clock_0/vdd clock_0/gnd clock_0/gnd clock_0/gnd clock_0/gnd clock_0/gnd
+ clock_0/vdd clock_0/gnd clock_0/gnd clock_0/vdd clock_0/vdd clock_0/gnd clock_0/vdd
+ clock_0/vdd clock_0/vdd clock_0/vdd clock_0/gnd clock_0/vdd clock_0/gnd clock_0/gnd
+ clock_0/gnd clock_0/gnd clock_0/gnd clock_0/vdd clock_0/vdd clock_0/vdd clock_0/vdd
+ clock_0/gnd clock_0/vdd clock_0/vdd clock_0/vdd clock_0/vdd clock_0/gnd clock_0/vdd
+ clock_0/gnd clock_0/vdd clock_0/vdd clock_0/gnd clock_0/gnd clock_0/vdd clock_0/gnd
+ clock_0/gnd clock_0/vdd clock_0/vdd clock_0/vdd clock_0/gnd clock_0/gnd clock_0/vdd
+ clock_0/gnd clock_0/gnd clock_0/gnd clock_0/vdd clock_0/vdd clock_0/gnd clock_0/vdd
+ clock_0/vdd clock_0/vdd clock_0/gnd clock_0/vdd clock_0/vdd clock_0/gnd clock_0/gnd
+ clock_0/gnd clock_0/vdd clock_0/vdd clock_0/vdd clock_0/gnd clock_0/vdd clock_0/vdd
+ clock_0/vdd clock_0/vdd clock_0/vdd clock_0/vdd clock_0/gnd clock_0/vdd clock_0/gnd
+ clock_0/vdd clock_0/gnd clock_0/gnd clock_0/gnd sky130_fd_pr__nfet_01v8_NJGC8F
Xsky130_fd_pr__nfet_01v8_NJGC8F_1 clock_0/vdd clock_0/gnd clock_0/gnd clock_0/vdd
+ clock_0/vdd clock_0/gnd clock_0/gnd clock_0/vdd clock_0/gnd clock_0/vdd clock_0/gnd
+ clock_0/gnd clock_0/vdd clock_0/gnd clock_0/gnd clock_0/gnd clock_0/vdd clock_0/gnd
+ clock_0/vdd clock_0/vdd clock_0/gnd clock_0/vdd clock_0/vdd clock_0/vdd clock_0/vdd
+ clock_0/gnd clock_0/vdd clock_0/vdd clock_0/gnd clock_0/vdd clock_0/vdd clock_0/gnd
+ clock_0/gnd clock_0/gnd clock_0/gnd clock_0/gnd clock_0/vdd clock_0/gnd clock_0/gnd
+ clock_0/vdd clock_0/gnd clock_0/gnd clock_0/gnd clock_0/vdd clock_0/gnd clock_0/gnd
+ clock_0/vdd clock_0/gnd clock_0/gnd clock_0/gnd clock_0/vdd clock_0/vdd clock_0/gnd
+ clock_0/gnd clock_0/vdd clock_0/gnd clock_0/gnd clock_0/vdd clock_0/gnd clock_0/gnd
+ clock_0/gnd clock_0/vdd clock_0/vdd clock_0/vdd clock_0/gnd clock_0/gnd clock_0/gnd
+ clock_0/gnd clock_0/vdd clock_0/gnd clock_0/vdd clock_0/gnd clock_0/vdd clock_0/gnd
+ clock_0/gnd clock_0/vdd clock_0/gnd clock_0/vdd clock_0/vdd clock_0/vdd clock_0/vdd
+ clock_0/vdd clock_0/vdd clock_0/gnd clock_0/gnd clock_0/gnd clock_0/gnd clock_0/gnd
+ clock_0/vdd clock_0/gnd clock_0/gnd clock_0/vdd clock_0/vdd clock_0/gnd clock_0/vdd
+ clock_0/vdd clock_0/vdd clock_0/vdd clock_0/gnd clock_0/vdd clock_0/gnd clock_0/gnd
+ clock_0/gnd clock_0/gnd clock_0/gnd clock_0/vdd clock_0/vdd clock_0/vdd clock_0/vdd
+ clock_0/gnd clock_0/vdd clock_0/vdd clock_0/vdd clock_0/vdd clock_0/gnd clock_0/vdd
+ clock_0/gnd clock_0/vdd clock_0/vdd clock_0/gnd clock_0/gnd clock_0/vdd clock_0/gnd
+ clock_0/gnd clock_0/vdd clock_0/vdd clock_0/vdd clock_0/gnd clock_0/gnd clock_0/vdd
+ clock_0/gnd clock_0/gnd clock_0/gnd clock_0/vdd clock_0/vdd clock_0/gnd clock_0/vdd
+ clock_0/vdd clock_0/vdd clock_0/gnd clock_0/vdd clock_0/vdd clock_0/gnd clock_0/gnd
+ clock_0/gnd clock_0/vdd clock_0/vdd clock_0/vdd clock_0/gnd clock_0/vdd clock_0/vdd
+ clock_0/vdd clock_0/vdd clock_0/vdd clock_0/vdd clock_0/gnd clock_0/vdd clock_0/gnd
+ clock_0/vdd clock_0/gnd clock_0/gnd clock_0/gnd sky130_fd_pr__nfet_01v8_NJGC8F
Xnmos_diode2_0 m1_12174_n760# nmos_dnw3_0/out2 nmos_dnw3_0/out1 nmos_dnw3_0/vs clock_0/gnd
+ nmos_diode2
Xsky130_fd_pr__cap_mim_m3_1_MH6KF8_0 nmos_dnw3_0/out2 clock_0/clkb clock_0/gnd sky130_fd_pr__cap_mim_m3_1_MH6KF8
Xsky130_fd_pr__cap_mim_m3_1_MH6KF8_1 nmos_dnw3_0/out1 clock_0/clk clock_0/gnd sky130_fd_pr__cap_mim_m3_1_MH6KF8
C0 nmos_dnw3_0/vs nmos_dnw3_0/out2 5.03f
C1 nmos_dnw3_0/out1 nmos_dnw3_0/out2 8.76f
C2 clock_0/vdd clock_0/clkb 18.1f
C3 nmos_dnw3_0/out1 nmos_dnw3_0/vs 3.18f
C4 clock_0/gnd clock_0/vdd 20.9f
C5 nmos_dnw3_0/vin clock_0/vdd 5.72f
C6 clock_0/clk clock_0/vdd 27.5f
C7 m1_12174_n760# clock_0/vdd 2.9f
C8 nmos_dnw3_0/vs 0 16.4f
C9 m1_12174_n760# 0 2.03f
C10 clock_0/a_2432_n962# 0 8.68f **FLOATING
C11 clock_0/a_2020_n482# 0 2.57f **FLOATING
C12 clock_0/a_344_102# 0 2.81f
C13 clock_0/a_2402_572# 0 2.17f
C14 clock_0/a_344_n986# 0 2.38f
C15 clock_0/a_3246_118# 0 6.83f
C16 nmos_dnw3_0/vin 0 2.2f
C17 nmos_dnw3_0/clkb 0 2.54f
C18 capacitors_5_0/capacitor_5_4/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C19 capacitors_5_0/capacitor_5_4/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C20 capacitors_5_0/capacitor_5_4/buffer_and_gate_0/in1 0 2.57f
C21 capacitors_5_0/capacitor_5_3/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C22 capacitors_5_0/capacitor_5_3/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C23 capacitors_5_0/capacitor_5_3/buffer_and_gate_0/in1 0 2.57f
C24 capacitors_5_0/capacitor_5_2/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C25 capacitors_5_0/capacitor_5_2/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C26 capacitors_5_0/capacitor_5_2/buffer_and_gate_0/in1 0 2.57f
C27 capacitors_5_0/capacitor_5_1/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C28 capacitors_5_0/capacitor_5_1/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C29 capacitors_5_0/capacitor_5_1/buffer_and_gate_0/in1 0 2.57f
C30 capacitors_5_0/capacitor_5_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C31 capacitors_5_0/capacitor_5_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C32 capacitors_5_0/capacitor_5_0/buffer_and_gate_0/in1 0 2.57f
C33 nmos_dnw3_0/out1 0 15f
C34 capacitors_5_0/capacitor_5_7/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C35 clock_0/clk 0 78.7f
C36 capacitors_5_0/capacitor_5_7/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C37 clock_0/gnd 0 0.12p
C38 capacitors_5_0/capacitor_5_7/buffer_and_gate_0/in1 0 2.57f
C39 capacitors_5_0/capacitor_5_6/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C40 capacitors_5_0/capacitor_5_6/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C41 capacitors_5_0/capacitor_5_6/buffer_and_gate_0/in1 0 2.57f
C42 capacitors_5_0/capacitor_5_5/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C43 capacitors_5_0/capacitor_5_5/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C44 capacitors_5_0/capacitor_5_5/buffer_and_gate_0/in1 0 2.57f
C45 capacitors_5_1/capacitor_5_4/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C46 capacitors_5_1/capacitor_5_4/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C47 capacitors_5_1/capacitor_5_4/buffer_and_gate_0/in1 0 2.57f
C48 capacitors_5_1/capacitor_5_3/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C49 capacitors_5_1/capacitor_5_3/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C50 capacitors_5_1/capacitor_5_3/buffer_and_gate_0/in1 0 2.57f
C51 capacitors_5_1/capacitor_5_2/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C52 capacitors_5_1/capacitor_5_2/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C53 capacitors_5_1/capacitor_5_2/buffer_and_gate_0/in1 0 2.57f
C54 capacitors_5_1/capacitor_5_1/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C55 capacitors_5_1/capacitor_5_1/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C56 capacitors_5_1/capacitor_5_1/buffer_and_gate_0/in1 0 2.57f
C57 capacitors_5_1/capacitor_5_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C58 capacitors_5_1/capacitor_5_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C59 capacitors_5_1/capacitor_5_0/buffer_and_gate_0/in1 0 2.57f
C60 nmos_dnw3_0/out2 0 13.6f
C61 capacitors_5_1/capacitor_5_7/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C62 clock_0/clkb 0 80.5f
C63 capacitors_5_1/capacitor_5_7/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C64 clock_0/vdd 0 0.481p
C65 capacitors_5_1/capacitor_5_7/buffer_and_gate_0/in1 0 2.57f
C66 capacitors_5_1/capacitor_5_6/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C67 capacitors_5_1/capacitor_5_6/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C68 capacitors_5_1/capacitor_5_6/buffer_and_gate_0/in1 0 2.57f
C69 capacitors_5_1/capacitor_5_5/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C70 capacitors_5_1/capacitor_5_5/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C71 capacitors_5_1/capacitor_5_5/buffer_and_gate_0/in1 0 2.57f
C72 nmos_dnw3_0/clk 0 2.76f
.ends

.subckt charge_pump_reverse nmos_dnw3_0/out2 m1_12174_n760# nmos_dnw3_0/vin clock_0/vdd
+ m2_10362_3360# m2_10308_13784# clock_0/clk clock_0/gnd m2_10400_5448# m2_10266_15868#
+ clock_0/clk_in m2_10426_9616# m2_10388_7530# m2_10336_11702# nmos_dnw3_0/vs m2_10436_1276#
Xsky130_fd_pr__cap_mim_m3_1_MH6KF8_4 nmos_dnw3_0/clk clock_0/clkb clock_0/gnd sky130_fd_pr__cap_mim_m3_1_MH6KF8
Xsky130_fd_pr__cap_mim_m3_1_MH6KF8_5 nmos_dnw3_0/clkb clock_0/clk clock_0/gnd sky130_fd_pr__cap_mim_m3_1_MH6KF8
Xcapacitors_5_1 nmos_dnw3_0/out2 clock_0/vdd clock_0/vdd clock_0/vdd m2_10400_5448#
+ m2_10266_15868# m2_10336_11702# m2_10388_7530# m2_10362_3360# m2_10426_9616# clock_0/clk
+ clock_0/vdd m2_10308_13784# m2_10436_1276# clock_0/gnd clock_0/vdd capacitors_5
Xcapacitors_5_0 nmos_dnw3_0/out1 clock_0/vdd clock_0/vdd clock_0/vdd m2_10400_5448#
+ m2_10266_15868# m2_10336_11702# m2_10388_7530# m2_10362_3360# m2_10426_9616# clock_0/clkb
+ clock_0/vdd m2_10308_13784# m2_10436_1276# clock_0/gnd clock_0/vdd capacitors_5
Xnmos_dnw3_0 nmos_dnw3_0/vin nmos_dnw3_0/out1 nmos_dnw3_0/out2 nmos_dnw3_0/clk nmos_dnw3_0/clkb
+ nmos_dnw3_0/vs clock_0/gnd nmos_dnw3
Xclock_0 clock_0/clk_in clock_0/vdd clock_0/gnd clock_0/clk clock_0/clkb clock
Xsky130_fd_pr__pfet_01v8_4RPJ49_0 clock_0/gnd clock_0/vdd clock_0/vdd clock_0/gnd
+ clock_0/gnd clock_0/vdd clock_0/vdd clock_0/vdd clock_0/gnd clock_0/vdd clock_0/gnd
+ clock_0/gnd clock_0/vdd clock_0/gnd clock_0/gnd clock_0/gnd clock_0/vdd clock_0/vdd
+ clock_0/vdd clock_0/vdd clock_0/gnd clock_0/vdd clock_0/gnd clock_0/gnd clock_0/gnd
+ clock_0/gnd clock_0/gnd clock_0/gnd clock_0/gnd clock_0/vdd clock_0/gnd clock_0/vdd
+ clock_0/gnd clock_0/gnd clock_0/vdd clock_0/gnd clock_0/gnd clock_0/vdd clock_0/vdd
+ clock_0/gnd clock_0/vdd clock_0/gnd clock_0/gnd clock_0/vdd clock_0/gnd clock_0/gnd
+ clock_0/vdd clock_0/vdd clock_0/gnd clock_0/gnd clock_0/vdd clock_0/vdd clock_0/vdd
+ clock_0/gnd clock_0/gnd clock_0/vdd clock_0/vdd clock_0/gnd clock_0/gnd clock_0/vdd
+ clock_0/vdd clock_0/gnd clock_0/vdd clock_0/gnd sky130_fd_pr__pfet_01v8_4RPJ49_0/w_n3905_n142#
+ clock_0/gnd clock_0/gnd clock_0/gnd clock_0/vdd clock_0/gnd clock_0/gnd clock_0/gnd
+ clock_0/vdd clock_0/vdd clock_0/gnd clock_0/gnd clock_0/vdd clock_0/vdd clock_0/gnd
+ clock_0/gnd clock_0/vdd clock_0/vdd clock_0/gnd clock_0/gnd clock_0/gnd clock_0/vdd
+ clock_0/vdd clock_0/vdd clock_0/vdd clock_0/vdd clock_0/vdd clock_0/vdd clock_0/vdd
+ clock_0/vdd clock_0/gnd clock_0/gnd clock_0/vdd clock_0/vdd clock_0/vdd clock_0/gnd
+ clock_0/vdd clock_0/vdd clock_0/vdd clock_0/vdd clock_0/vdd clock_0/gnd clock_0/vdd
+ clock_0/vdd clock_0/gnd clock_0/vdd clock_0/vdd clock_0/gnd clock_0/gnd clock_0/gnd
+ clock_0/gnd clock_0/gnd clock_0/vdd clock_0/vdd clock_0/vdd clock_0/gnd clock_0/vdd
+ clock_0/vdd clock_0/gnd clock_0/vdd clock_0/gnd clock_0/vdd clock_0/vdd clock_0/vdd
+ clock_0/gnd clock_0/gnd clock_0/vdd clock_0/vdd clock_0/gnd clock_0/vdd clock_0/vdd
+ clock_0/vdd clock_0/vdd clock_0/gnd clock_0/vdd clock_0/gnd clock_0/gnd clock_0/gnd
+ clock_0/vdd clock_0/vdd clock_0/vdd clock_0/gnd clock_0/gnd clock_0/gnd clock_0/gnd
+ clock_0/vdd clock_0/gnd clock_0/gnd clock_0/gnd clock_0/vdd clock_0/gnd clock_0/gnd
+ clock_0/gnd clock_0/gnd clock_0/vdd clock_0/gnd clock_0/gnd clock_0/vdd clock_0/vdd
+ sky130_fd_pr__pfet_01v8_4RPJ49
Xsky130_fd_pr__pfet_01v8_4RPJ49_1 clock_0/gnd clock_0/vdd clock_0/vdd clock_0/gnd
+ clock_0/gnd clock_0/vdd clock_0/vdd clock_0/vdd clock_0/gnd clock_0/vdd clock_0/gnd
+ clock_0/gnd clock_0/vdd clock_0/gnd clock_0/gnd clock_0/gnd clock_0/vdd clock_0/vdd
+ clock_0/vdd clock_0/vdd clock_0/gnd clock_0/vdd clock_0/gnd clock_0/gnd clock_0/gnd
+ clock_0/gnd clock_0/gnd clock_0/gnd clock_0/gnd clock_0/vdd clock_0/gnd clock_0/vdd
+ clock_0/gnd clock_0/gnd clock_0/vdd clock_0/gnd clock_0/gnd clock_0/vdd clock_0/vdd
+ clock_0/gnd clock_0/vdd clock_0/gnd clock_0/gnd clock_0/vdd clock_0/gnd clock_0/gnd
+ clock_0/vdd clock_0/vdd clock_0/gnd clock_0/gnd clock_0/vdd clock_0/vdd clock_0/vdd
+ clock_0/gnd clock_0/gnd clock_0/vdd clock_0/vdd clock_0/gnd clock_0/gnd clock_0/vdd
+ clock_0/vdd clock_0/gnd clock_0/vdd clock_0/gnd sky130_fd_pr__pfet_01v8_4RPJ49_1/w_n3905_n142#
+ clock_0/gnd clock_0/gnd clock_0/gnd clock_0/vdd clock_0/gnd clock_0/gnd clock_0/gnd
+ clock_0/vdd clock_0/vdd clock_0/gnd clock_0/gnd clock_0/vdd clock_0/vdd clock_0/gnd
+ clock_0/gnd clock_0/vdd clock_0/vdd clock_0/gnd clock_0/gnd clock_0/gnd clock_0/vdd
+ clock_0/vdd clock_0/vdd clock_0/vdd clock_0/vdd clock_0/vdd clock_0/vdd clock_0/vdd
+ clock_0/vdd clock_0/gnd clock_0/gnd clock_0/vdd clock_0/vdd clock_0/vdd clock_0/gnd
+ clock_0/vdd clock_0/vdd clock_0/vdd clock_0/vdd clock_0/vdd clock_0/gnd clock_0/vdd
+ clock_0/vdd clock_0/gnd clock_0/vdd clock_0/vdd clock_0/gnd clock_0/gnd clock_0/gnd
+ clock_0/gnd clock_0/gnd clock_0/vdd clock_0/vdd clock_0/vdd clock_0/gnd clock_0/vdd
+ clock_0/vdd clock_0/gnd clock_0/vdd clock_0/gnd clock_0/vdd clock_0/vdd clock_0/vdd
+ clock_0/gnd clock_0/gnd clock_0/vdd clock_0/vdd clock_0/gnd clock_0/vdd clock_0/vdd
+ clock_0/vdd clock_0/vdd clock_0/gnd clock_0/vdd clock_0/gnd clock_0/gnd clock_0/gnd
+ clock_0/vdd clock_0/vdd clock_0/vdd clock_0/gnd clock_0/gnd clock_0/gnd clock_0/gnd
+ clock_0/vdd clock_0/gnd clock_0/gnd clock_0/gnd clock_0/vdd clock_0/gnd clock_0/gnd
+ clock_0/gnd clock_0/gnd clock_0/vdd clock_0/gnd clock_0/gnd clock_0/vdd clock_0/vdd
+ sky130_fd_pr__pfet_01v8_4RPJ49
Xsky130_fd_pr__nfet_01v8_NJGC8F_0 clock_0/vdd clock_0/gnd clock_0/gnd clock_0/vdd
+ clock_0/vdd clock_0/gnd clock_0/gnd clock_0/vdd clock_0/gnd clock_0/vdd clock_0/gnd
+ clock_0/gnd clock_0/vdd clock_0/gnd clock_0/gnd clock_0/gnd clock_0/vdd clock_0/gnd
+ clock_0/vdd clock_0/vdd clock_0/gnd clock_0/vdd clock_0/vdd clock_0/vdd clock_0/vdd
+ clock_0/gnd clock_0/vdd clock_0/vdd clock_0/gnd clock_0/vdd clock_0/vdd clock_0/gnd
+ clock_0/gnd clock_0/gnd clock_0/gnd clock_0/gnd clock_0/vdd clock_0/gnd clock_0/gnd
+ clock_0/vdd clock_0/gnd clock_0/gnd clock_0/gnd clock_0/vdd clock_0/gnd clock_0/gnd
+ clock_0/vdd clock_0/gnd clock_0/gnd clock_0/gnd clock_0/vdd clock_0/vdd clock_0/gnd
+ clock_0/gnd clock_0/vdd clock_0/gnd clock_0/gnd clock_0/vdd clock_0/gnd clock_0/gnd
+ clock_0/gnd clock_0/vdd clock_0/vdd clock_0/vdd clock_0/gnd clock_0/gnd clock_0/gnd
+ clock_0/gnd clock_0/vdd clock_0/gnd clock_0/vdd clock_0/gnd clock_0/vdd clock_0/gnd
+ clock_0/gnd clock_0/vdd clock_0/gnd clock_0/vdd clock_0/vdd clock_0/vdd clock_0/vdd
+ clock_0/vdd clock_0/vdd clock_0/gnd clock_0/gnd clock_0/gnd clock_0/gnd clock_0/gnd
+ clock_0/vdd clock_0/gnd clock_0/gnd clock_0/vdd clock_0/vdd clock_0/gnd clock_0/vdd
+ clock_0/vdd clock_0/vdd clock_0/vdd clock_0/gnd clock_0/vdd clock_0/gnd clock_0/gnd
+ clock_0/gnd clock_0/gnd clock_0/gnd clock_0/vdd clock_0/vdd clock_0/vdd clock_0/vdd
+ clock_0/gnd clock_0/vdd clock_0/vdd clock_0/vdd clock_0/vdd clock_0/gnd clock_0/vdd
+ clock_0/gnd clock_0/vdd clock_0/vdd clock_0/gnd clock_0/gnd clock_0/vdd clock_0/gnd
+ clock_0/gnd clock_0/vdd clock_0/vdd clock_0/vdd clock_0/gnd clock_0/gnd clock_0/vdd
+ clock_0/gnd clock_0/gnd clock_0/gnd clock_0/vdd clock_0/vdd clock_0/gnd clock_0/vdd
+ clock_0/vdd clock_0/vdd clock_0/gnd clock_0/vdd clock_0/vdd clock_0/gnd clock_0/gnd
+ clock_0/gnd clock_0/vdd clock_0/vdd clock_0/vdd clock_0/gnd clock_0/vdd clock_0/vdd
+ clock_0/vdd clock_0/vdd clock_0/vdd clock_0/vdd clock_0/gnd clock_0/vdd clock_0/gnd
+ clock_0/vdd clock_0/gnd clock_0/gnd clock_0/gnd sky130_fd_pr__nfet_01v8_NJGC8F
Xsky130_fd_pr__nfet_01v8_NJGC8F_1 clock_0/vdd clock_0/gnd clock_0/gnd clock_0/vdd
+ clock_0/vdd clock_0/gnd clock_0/gnd clock_0/vdd clock_0/gnd clock_0/vdd clock_0/gnd
+ clock_0/gnd clock_0/vdd clock_0/gnd clock_0/gnd clock_0/gnd clock_0/vdd clock_0/gnd
+ clock_0/vdd clock_0/vdd clock_0/gnd clock_0/vdd clock_0/vdd clock_0/vdd clock_0/vdd
+ clock_0/gnd clock_0/vdd clock_0/vdd clock_0/gnd clock_0/vdd clock_0/vdd clock_0/gnd
+ clock_0/gnd clock_0/gnd clock_0/gnd clock_0/gnd clock_0/vdd clock_0/gnd clock_0/gnd
+ clock_0/vdd clock_0/gnd clock_0/gnd clock_0/gnd clock_0/vdd clock_0/gnd clock_0/gnd
+ clock_0/vdd clock_0/gnd clock_0/gnd clock_0/gnd clock_0/vdd clock_0/vdd clock_0/gnd
+ clock_0/gnd clock_0/vdd clock_0/gnd clock_0/gnd clock_0/vdd clock_0/gnd clock_0/gnd
+ clock_0/gnd clock_0/vdd clock_0/vdd clock_0/vdd clock_0/gnd clock_0/gnd clock_0/gnd
+ clock_0/gnd clock_0/vdd clock_0/gnd clock_0/vdd clock_0/gnd clock_0/vdd clock_0/gnd
+ clock_0/gnd clock_0/vdd clock_0/gnd clock_0/vdd clock_0/vdd clock_0/vdd clock_0/vdd
+ clock_0/vdd clock_0/vdd clock_0/gnd clock_0/gnd clock_0/gnd clock_0/gnd clock_0/gnd
+ clock_0/vdd clock_0/gnd clock_0/gnd clock_0/vdd clock_0/vdd clock_0/gnd clock_0/vdd
+ clock_0/vdd clock_0/vdd clock_0/vdd clock_0/gnd clock_0/vdd clock_0/gnd clock_0/gnd
+ clock_0/gnd clock_0/gnd clock_0/gnd clock_0/vdd clock_0/vdd clock_0/vdd clock_0/vdd
+ clock_0/gnd clock_0/vdd clock_0/vdd clock_0/vdd clock_0/vdd clock_0/gnd clock_0/vdd
+ clock_0/gnd clock_0/vdd clock_0/vdd clock_0/gnd clock_0/gnd clock_0/vdd clock_0/gnd
+ clock_0/gnd clock_0/vdd clock_0/vdd clock_0/vdd clock_0/gnd clock_0/gnd clock_0/vdd
+ clock_0/gnd clock_0/gnd clock_0/gnd clock_0/vdd clock_0/vdd clock_0/gnd clock_0/vdd
+ clock_0/vdd clock_0/vdd clock_0/gnd clock_0/vdd clock_0/vdd clock_0/gnd clock_0/gnd
+ clock_0/gnd clock_0/vdd clock_0/vdd clock_0/vdd clock_0/gnd clock_0/vdd clock_0/vdd
+ clock_0/vdd clock_0/vdd clock_0/vdd clock_0/vdd clock_0/gnd clock_0/vdd clock_0/gnd
+ clock_0/vdd clock_0/gnd clock_0/gnd clock_0/gnd sky130_fd_pr__nfet_01v8_NJGC8F
Xnmos_diode2_0 m1_12174_n760# nmos_dnw3_0/out2 nmos_dnw3_0/out1 nmos_dnw3_0/vs clock_0/gnd
+ nmos_diode2
Xsky130_fd_pr__cap_mim_m3_1_MH6KF8_0 nmos_dnw3_0/out2 clock_0/clk clock_0/gnd sky130_fd_pr__cap_mim_m3_1_MH6KF8
Xsky130_fd_pr__cap_mim_m3_1_MH6KF8_1 nmos_dnw3_0/out1 clock_0/clkb clock_0/gnd sky130_fd_pr__cap_mim_m3_1_MH6KF8
C0 nmos_dnw3_0/vin clock_0/vdd 8.87f
C1 clock_0/clkb clock_0/vdd 24.4f
C2 nmos_dnw3_0/out1 nmos_dnw3_0/vs 3.18f
C3 m1_12174_n760# clock_0/vdd 2.66f
C4 nmos_dnw3_0/out2 nmos_dnw3_0/vs 5.03f
C5 nmos_dnw3_0/out1 nmos_dnw3_0/out2 8.76f
C6 clock_0/gnd clock_0/vdd 18.8f
C7 clock_0/clk clock_0/vdd 20f
C8 nmos_dnw3_0/vs 0 16.4f
C9 m1_12174_n760# 0 2.31f
C10 sky130_fd_pr__pfet_01v8_4RPJ49_1/w_n3905_n142# 0 6.63f
C11 sky130_fd_pr__pfet_01v8_4RPJ49_0/w_n3905_n142# 0 6.63f
C12 clock_0/a_2432_n962# 0 8.68f **FLOATING
C13 clock_0/a_2020_n482# 0 2.57f **FLOATING
C14 clock_0/a_344_102# 0 2.81f
C15 clock_0/a_2402_572# 0 2.17f
C16 clock_0/a_344_n986# 0 2.38f
C17 clock_0/a_3246_118# 0 6.83f
C18 nmos_dnw3_0/vin 0 2.47f
C19 nmos_dnw3_0/clkb 0 2.23f
C20 capacitors_5_0/capacitor_5_4/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C21 capacitors_5_0/capacitor_5_4/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C22 capacitors_5_0/capacitor_5_4/buffer_and_gate_0/in1 0 2.57f
C23 capacitors_5_0/capacitor_5_3/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C24 capacitors_5_0/capacitor_5_3/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C25 capacitors_5_0/capacitor_5_3/buffer_and_gate_0/in1 0 2.57f
C26 capacitors_5_0/capacitor_5_2/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C27 capacitors_5_0/capacitor_5_2/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C28 capacitors_5_0/capacitor_5_2/buffer_and_gate_0/in1 0 2.57f
C29 capacitors_5_0/capacitor_5_1/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C30 capacitors_5_0/capacitor_5_1/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C31 capacitors_5_0/capacitor_5_1/buffer_and_gate_0/in1 0 2.57f
C32 capacitors_5_0/capacitor_5_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C33 capacitors_5_0/capacitor_5_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C34 capacitors_5_0/capacitor_5_0/buffer_and_gate_0/in1 0 2.57f
C35 nmos_dnw3_0/out1 0 15.1f
C36 capacitors_5_0/capacitor_5_7/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C37 clock_0/clkb 0 86.4f
C38 capacitors_5_0/capacitor_5_7/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C39 capacitors_5_0/capacitor_5_7/buffer_and_gate_0/in1 0 2.57f
C40 capacitors_5_0/capacitor_5_6/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C41 capacitors_5_0/capacitor_5_6/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C42 capacitors_5_0/capacitor_5_6/buffer_and_gate_0/in1 0 2.57f
C43 capacitors_5_0/capacitor_5_5/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C44 capacitors_5_0/capacitor_5_5/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C45 capacitors_5_0/capacitor_5_5/buffer_and_gate_0/in1 0 2.57f
C46 capacitors_5_1/capacitor_5_4/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C47 capacitors_5_1/capacitor_5_4/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C48 capacitors_5_1/capacitor_5_4/buffer_and_gate_0/in1 0 2.57f
C49 capacitors_5_1/capacitor_5_3/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C50 capacitors_5_1/capacitor_5_3/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C51 capacitors_5_1/capacitor_5_3/buffer_and_gate_0/in1 0 2.57f
C52 capacitors_5_1/capacitor_5_2/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C53 capacitors_5_1/capacitor_5_2/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C54 capacitors_5_1/capacitor_5_2/buffer_and_gate_0/in1 0 2.57f
C55 capacitors_5_1/capacitor_5_1/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C56 capacitors_5_1/capacitor_5_1/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C57 capacitors_5_1/capacitor_5_1/buffer_and_gate_0/in1 0 2.57f
C58 capacitors_5_1/capacitor_5_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C59 capacitors_5_1/capacitor_5_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C60 capacitors_5_1/capacitor_5_0/buffer_and_gate_0/in1 0 2.57f
C61 nmos_dnw3_0/out2 0 14.9f
C62 capacitors_5_1/capacitor_5_7/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C63 clock_0/clk 0 80f
C64 capacitors_5_1/capacitor_5_7/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C65 clock_0/vdd 0 0.466p
C66 clock_0/gnd 0 0.116p
C67 capacitors_5_1/capacitor_5_7/buffer_and_gate_0/in1 0 2.57f
C68 capacitors_5_1/capacitor_5_6/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C69 capacitors_5_1/capacitor_5_6/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C70 capacitors_5_1/capacitor_5_6/buffer_and_gate_0/in1 0 2.57f
C71 capacitors_5_1/capacitor_5_5/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C72 capacitors_5_1/capacitor_5_5/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C73 capacitors_5_1/capacitor_5_5/buffer_and_gate_0/in1 0 2.57f
C74 nmos_dnw3_0/clk 0 2.43f
.ends

.subckt CP2_5_stage charge_pump_reverse_1/nmos_dnw3_0/vs m1_94493_n2143# charge_pump_reverse_1/nmos_dnw3_0/out2
+ m1_71529_n2069# charge_pump_2/m1_12174_n760# charge_pump_reverse_0/nmos_dnw3_0/vin
+ charge_pump_2/clock_0/vdd m2_91760_11118# charge_pump_0/nmos_dnw3_0/vin m2_91682_21576#
+ charge_pump_0/nmos_dnw3_0/vs charge_pump_reverse_1/clock_0/clk m2_91774_13212# m2_91694_23658#
+ charge_pump_2/nmos_dnw3_0/vs m2_91690_17386# charge_pump_1/nmos_dnw3_0/vs charge_pump_reverse_0/nmos_dnw3_0/vs
+ m2_91686_15288# charge_pump_2/clock_0/clk_in charge_pump_0/clock_0/clk_in charge_pump_reverse_1/clock_0/clk_in
+ m2_91764_9020# m2_91690_19482# VSUBS
Xcharge_pump_0 charge_pump_reverse_0/nmos_dnw3_0/vin charge_pump_0/nmos_dnw3_0/vin
+ m2_91690_17386# charge_pump_0/clock_0/clk_in m2_91774_13212# m2_91686_15288# m2_91694_23658#
+ m2_91690_19482# m2_91764_9020# m2_91760_11118# m2_91682_21576# charge_pump_2/clock_0/vdd
+ charge_pump_0/nmos_dnw3_0/vs VSUBS charge_pump
Xcharge_pump_1 charge_pump_reverse_1/nmos_dnw3_0/vin charge_pump_1/nmos_dnw3_0/vin
+ m2_91690_17386# charge_pump_1/clock_0/clk_in m2_91774_13212# m2_91686_15288# m2_91694_23658#
+ m2_91690_19482# m2_91764_9020# m2_91760_11118# m2_91682_21576# charge_pump_2/clock_0/vdd
+ charge_pump_1/nmos_dnw3_0/vs VSUBS charge_pump
Xbuffer_digital_0 m1_20940_n2218# buffer_digital_0/a_116_148# charge_pump_2/clock_0/vdd
+ charge_pump_2/clock_0/vdd charge_pump_0/clock_0/clk_in VSUBS VSUBS VSUBS buffer_digital
Xcharge_pump_2 charge_pump_2/m1_12174_n760# charge_pump_2/nmos_dnw3_0/vin m2_91690_17386#
+ charge_pump_2/clock_0/clk_in m2_91774_13212# m2_91686_15288# m2_91694_23658# m2_91690_19482#
+ m2_91764_9020# m2_91760_11118# m2_91682_21576# charge_pump_2/clock_0/vdd charge_pump_2/nmos_dnw3_0/vs
+ VSUBS charge_pump
Xbuffer_digital_1 charge_pump_reverse_0/clock_0/clk_in buffer_digital_1/a_116_148#
+ charge_pump_2/clock_0/vdd charge_pump_2/clock_0/vdd m1_20940_n2218# VSUBS VSUBS
+ VSUBS buffer_digital
Xbuffer_digital_2 m1_45014_n2098# buffer_digital_2/a_116_148# charge_pump_2/clock_0/vdd
+ charge_pump_2/clock_0/vdd charge_pump_reverse_0/clock_0/clk_in VSUBS VSUBS VSUBS
+ buffer_digital
Xbuffer_digital_3 charge_pump_1/clock_0/clk_in buffer_digital_3/a_116_148# charge_pump_2/clock_0/vdd
+ charge_pump_2/clock_0/vdd m1_45014_n2098# VSUBS VSUBS VSUBS buffer_digital
Xbuffer_digital_5 m1_71529_n2069# buffer_digital_5/a_116_148# charge_pump_2/clock_0/vdd
+ charge_pump_2/clock_0/vdd m1_68586_n2076# buffer_digital_5/m1_n2_0# buffer_digital_5/m1_216_0#
+ VSUBS buffer_digital
Xbuffer_digital_4 m1_68586_n2076# buffer_digital_4/a_116_148# charge_pump_2/clock_0/vdd
+ charge_pump_2/clock_0/vdd charge_pump_1/clock_0/clk_in VSUBS buffer_digital_4/m1_216_0#
+ VSUBS buffer_digital
Xbuffer_digital_6 m1_91387_n2165# buffer_digital_6/a_116_148# charge_pump_2/clock_0/vdd
+ charge_pump_2/clock_0/vdd m1_71529_n2069# VSUBS VSUBS VSUBS buffer_digital
Xbuffer_digital_7 m1_94493_n2143# buffer_digital_7/a_116_148# charge_pump_2/clock_0/vdd
+ charge_pump_2/clock_0/vdd m1_91387_n2165# VSUBS VSUBS VSUBS buffer_digital
Xcharge_pump_reverse_0 charge_pump_reverse_0/nmos_dnw3_0/out2 charge_pump_1/nmos_dnw3_0/vin
+ charge_pump_reverse_0/nmos_dnw3_0/vin charge_pump_2/clock_0/vdd m2_91682_21576#
+ m2_91760_11118# charge_pump_reverse_0/clock_0/clk VSUBS m2_91690_19482# m2_91764_9020#
+ charge_pump_reverse_0/clock_0/clk_in m2_91686_15288# m2_91690_17386# m2_91774_13212#
+ charge_pump_reverse_0/nmos_dnw3_0/vs m2_91694_23658# charge_pump_reverse
Xcharge_pump_reverse_1 charge_pump_reverse_1/nmos_dnw3_0/out2 charge_pump_2/nmos_dnw3_0/vin
+ charge_pump_reverse_1/nmos_dnw3_0/vin charge_pump_2/clock_0/vdd m2_91682_21576#
+ m2_91760_11118# charge_pump_reverse_1/clock_0/clk VSUBS m2_91690_19482# m2_91764_9020#
+ charge_pump_reverse_1/clock_0/clk_in m2_91686_15288# m2_91690_17386# m2_91774_13212#
+ charge_pump_reverse_1/nmos_dnw3_0/vs m2_91694_23658# charge_pump_reverse
C0 charge_pump_2/clock_0/vdd m2_91764_9020# 4.32f
C1 charge_pump_2/clock_0/vdd m2_91682_21576# 4.18f
C2 m2_91760_11118# VSUBS 4.15f
C3 VSUBS m2_91694_23658# 3f
C4 VSUBS m2_91686_15288# 4.14f
C5 VSUBS m2_91690_19482# 4.16f
C6 m2_91774_13212# VSUBS 4.04f
C7 charge_pump_2/clock_0/vdd charge_pump_0/clock_0/clk_in 4.51f
C8 m2_91760_11118# charge_pump_2/clock_0/vdd 4.28f
C9 charge_pump_2/clock_0/vdd charge_pump_1/clock_0/clk_in 4.25f
C10 charge_pump_2/clock_0/vdd m2_91694_23658# 4.11f
C11 charge_pump_2/clock_0/vdd m2_91686_15288# 4.26f
C12 VSUBS m2_91690_17386# 4.15f
C13 charge_pump_2/clock_0/vdd m1_71529_n2069# 4.34f
C14 charge_pump_2/clock_0/vdd m2_91690_19482# 4.29f
C15 charge_pump_2/clock_0/vdd charge_pump_reverse_0/clock_0/clk_in 4.33f
C16 m2_91774_13212# charge_pump_2/clock_0/vdd 4.17f
C17 charge_pump_2/clock_0/vdd m1_94493_n2143# 2.17f
C18 VSUBS m2_91764_9020# 3.2f
C19 charge_pump_2/clock_0/vdd m2_91690_17386# 4.27f
C20 charge_pump_2/clock_0/vdd VSUBS 26.7f
C21 VSUBS m2_91682_21576# 4.04f
C22 charge_pump_reverse_1/nmos_dnw3_0/vs 0 16.4f
C23 charge_pump_reverse_1/sky130_fd_pr__pfet_01v8_4RPJ49_1/w_n3905_n142# 0 6.63f
C24 charge_pump_reverse_1/sky130_fd_pr__pfet_01v8_4RPJ49_0/w_n3905_n142# 0 6.63f
C25 charge_pump_reverse_1/clock_0/a_2432_n962# 0 8.68f **FLOATING
C26 charge_pump_reverse_1/clock_0/a_2020_n482# 0 2.57f **FLOATING
C27 charge_pump_reverse_1/clock_0/a_344_102# 0 2.81f
C28 charge_pump_reverse_1/clock_0/a_2402_572# 0 2.17f
C29 charge_pump_reverse_1/clock_0/a_344_n986# 0 2.38f
C30 charge_pump_reverse_1/clock_0/a_3246_118# 0 6.83f
C31 charge_pump_reverse_1/nmos_dnw3_0/clkb 0 2.23f
C32 charge_pump_reverse_1/capacitors_5_0/capacitor_5_4/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C33 charge_pump_reverse_1/capacitors_5_0/capacitor_5_4/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C34 charge_pump_reverse_1/capacitors_5_0/capacitor_5_4/buffer_and_gate_0/in1 0 2.57f
C35 charge_pump_reverse_1/capacitors_5_0/capacitor_5_3/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C36 charge_pump_reverse_1/capacitors_5_0/capacitor_5_3/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C37 charge_pump_reverse_1/capacitors_5_0/capacitor_5_3/buffer_and_gate_0/in1 0 2.57f
C38 charge_pump_reverse_1/capacitors_5_0/capacitor_5_2/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C39 charge_pump_reverse_1/capacitors_5_0/capacitor_5_2/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C40 charge_pump_reverse_1/capacitors_5_0/capacitor_5_2/buffer_and_gate_0/in1 0 2.57f
C41 charge_pump_reverse_1/capacitors_5_0/capacitor_5_1/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C42 charge_pump_reverse_1/capacitors_5_0/capacitor_5_1/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C43 charge_pump_reverse_1/capacitors_5_0/capacitor_5_1/buffer_and_gate_0/in1 0 2.57f
C44 charge_pump_reverse_1/capacitors_5_0/capacitor_5_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C45 charge_pump_reverse_1/capacitors_5_0/capacitor_5_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C46 charge_pump_reverse_1/capacitors_5_0/capacitor_5_0/buffer_and_gate_0/in1 0 2.57f
C47 charge_pump_reverse_1/nmos_dnw3_0/out1 0 15.1f
C48 charge_pump_reverse_1/capacitors_5_0/capacitor_5_7/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C49 charge_pump_reverse_1/clock_0/clkb 0 86.4f
C50 charge_pump_reverse_1/capacitors_5_0/capacitor_5_7/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C51 charge_pump_reverse_1/capacitors_5_0/capacitor_5_7/buffer_and_gate_0/in1 0 2.57f
C52 charge_pump_reverse_1/capacitors_5_0/capacitor_5_6/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C53 charge_pump_reverse_1/capacitors_5_0/capacitor_5_6/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C54 charge_pump_reverse_1/capacitors_5_0/capacitor_5_6/buffer_and_gate_0/in1 0 2.57f
C55 charge_pump_reverse_1/capacitors_5_0/capacitor_5_5/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C56 charge_pump_reverse_1/capacitors_5_0/capacitor_5_5/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C57 charge_pump_reverse_1/capacitors_5_0/capacitor_5_5/buffer_and_gate_0/in1 0 2.57f
C58 charge_pump_reverse_1/capacitors_5_1/capacitor_5_4/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C59 charge_pump_reverse_1/capacitors_5_1/capacitor_5_4/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C60 charge_pump_reverse_1/capacitors_5_1/capacitor_5_4/buffer_and_gate_0/in1 0 2.57f
C61 charge_pump_reverse_1/capacitors_5_1/capacitor_5_3/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C62 charge_pump_reverse_1/capacitors_5_1/capacitor_5_3/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C63 charge_pump_reverse_1/capacitors_5_1/capacitor_5_3/buffer_and_gate_0/in1 0 2.57f
C64 charge_pump_reverse_1/capacitors_5_1/capacitor_5_2/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C65 charge_pump_reverse_1/capacitors_5_1/capacitor_5_2/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C66 charge_pump_reverse_1/capacitors_5_1/capacitor_5_2/buffer_and_gate_0/in1 0 2.57f
C67 charge_pump_reverse_1/capacitors_5_1/capacitor_5_1/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C68 charge_pump_reverse_1/capacitors_5_1/capacitor_5_1/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C69 charge_pump_reverse_1/capacitors_5_1/capacitor_5_1/buffer_and_gate_0/in1 0 2.57f
C70 charge_pump_reverse_1/capacitors_5_1/capacitor_5_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C71 charge_pump_reverse_1/capacitors_5_1/capacitor_5_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C72 charge_pump_reverse_1/capacitors_5_1/capacitor_5_0/buffer_and_gate_0/in1 0 2.57f
C73 charge_pump_reverse_1/nmos_dnw3_0/out2 0 14.9f
C74 charge_pump_reverse_1/capacitors_5_1/capacitor_5_7/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C75 charge_pump_reverse_1/clock_0/clk 0 80f
C76 charge_pump_reverse_1/capacitors_5_1/capacitor_5_7/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C77 charge_pump_reverse_1/capacitors_5_1/capacitor_5_7/buffer_and_gate_0/in1 0 2.57f
C78 charge_pump_reverse_1/capacitors_5_1/capacitor_5_6/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C79 charge_pump_reverse_1/capacitors_5_1/capacitor_5_6/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C80 charge_pump_reverse_1/capacitors_5_1/capacitor_5_6/buffer_and_gate_0/in1 0 2.57f
C81 charge_pump_reverse_1/capacitors_5_1/capacitor_5_5/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C82 charge_pump_reverse_1/capacitors_5_1/capacitor_5_5/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C83 charge_pump_reverse_1/capacitors_5_1/capacitor_5_5/buffer_and_gate_0/in1 0 2.57f
C84 charge_pump_reverse_1/nmos_dnw3_0/clk 0 2.43f
C85 charge_pump_reverse_0/nmos_dnw3_0/vs 0 16.4f
C86 charge_pump_reverse_0/sky130_fd_pr__pfet_01v8_4RPJ49_1/w_n3905_n142# 0 6.63f
C87 charge_pump_reverse_0/sky130_fd_pr__pfet_01v8_4RPJ49_0/w_n3905_n142# 0 6.63f
C88 charge_pump_reverse_0/clock_0/a_2432_n962# 0 8.68f **FLOATING
C89 charge_pump_reverse_0/clock_0/a_2020_n482# 0 2.57f **FLOATING
C90 charge_pump_reverse_0/clock_0/a_344_102# 0 2.81f
C91 charge_pump_reverse_0/clock_0/a_2402_572# 0 2.17f
C92 charge_pump_reverse_0/clock_0/a_344_n986# 0 2.38f
C93 charge_pump_reverse_0/clock_0/a_3246_118# 0 6.83f
C94 charge_pump_reverse_0/nmos_dnw3_0/clkb 0 2.23f
C95 charge_pump_reverse_0/capacitors_5_0/capacitor_5_4/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C96 charge_pump_reverse_0/capacitors_5_0/capacitor_5_4/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C97 charge_pump_reverse_0/capacitors_5_0/capacitor_5_4/buffer_and_gate_0/in1 0 2.57f
C98 charge_pump_reverse_0/capacitors_5_0/capacitor_5_3/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C99 charge_pump_reverse_0/capacitors_5_0/capacitor_5_3/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C100 charge_pump_reverse_0/capacitors_5_0/capacitor_5_3/buffer_and_gate_0/in1 0 2.57f
C101 charge_pump_reverse_0/capacitors_5_0/capacitor_5_2/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C102 charge_pump_reverse_0/capacitors_5_0/capacitor_5_2/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C103 charge_pump_reverse_0/capacitors_5_0/capacitor_5_2/buffer_and_gate_0/in1 0 2.57f
C104 charge_pump_reverse_0/capacitors_5_0/capacitor_5_1/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C105 charge_pump_reverse_0/capacitors_5_0/capacitor_5_1/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C106 charge_pump_reverse_0/capacitors_5_0/capacitor_5_1/buffer_and_gate_0/in1 0 2.57f
C107 charge_pump_reverse_0/capacitors_5_0/capacitor_5_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C108 charge_pump_reverse_0/capacitors_5_0/capacitor_5_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C109 charge_pump_reverse_0/capacitors_5_0/capacitor_5_0/buffer_and_gate_0/in1 0 2.57f
C110 charge_pump_reverse_0/nmos_dnw3_0/out1 0 15.1f
C111 charge_pump_reverse_0/capacitors_5_0/capacitor_5_7/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C112 charge_pump_reverse_0/clock_0/clkb 0 86.4f
C113 charge_pump_reverse_0/capacitors_5_0/capacitor_5_7/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C114 charge_pump_reverse_0/capacitors_5_0/capacitor_5_7/buffer_and_gate_0/in1 0 2.57f
C115 charge_pump_reverse_0/capacitors_5_0/capacitor_5_6/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C116 charge_pump_reverse_0/capacitors_5_0/capacitor_5_6/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C117 charge_pump_reverse_0/capacitors_5_0/capacitor_5_6/buffer_and_gate_0/in1 0 2.57f
C118 charge_pump_reverse_0/capacitors_5_0/capacitor_5_5/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C119 charge_pump_reverse_0/capacitors_5_0/capacitor_5_5/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C120 charge_pump_reverse_0/capacitors_5_0/capacitor_5_5/buffer_and_gate_0/in1 0 2.57f
C121 charge_pump_reverse_0/capacitors_5_1/capacitor_5_4/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C122 charge_pump_reverse_0/capacitors_5_1/capacitor_5_4/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C123 charge_pump_reverse_0/capacitors_5_1/capacitor_5_4/buffer_and_gate_0/in1 0 2.57f
C124 charge_pump_reverse_0/capacitors_5_1/capacitor_5_3/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C125 charge_pump_reverse_0/capacitors_5_1/capacitor_5_3/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C126 charge_pump_reverse_0/capacitors_5_1/capacitor_5_3/buffer_and_gate_0/in1 0 2.57f
C127 charge_pump_reverse_0/capacitors_5_1/capacitor_5_2/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C128 charge_pump_reverse_0/capacitors_5_1/capacitor_5_2/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C129 charge_pump_reverse_0/capacitors_5_1/capacitor_5_2/buffer_and_gate_0/in1 0 2.57f
C130 charge_pump_reverse_0/capacitors_5_1/capacitor_5_1/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C131 charge_pump_reverse_0/capacitors_5_1/capacitor_5_1/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C132 charge_pump_reverse_0/capacitors_5_1/capacitor_5_1/buffer_and_gate_0/in1 0 2.57f
C133 charge_pump_reverse_0/capacitors_5_1/capacitor_5_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C134 charge_pump_reverse_0/capacitors_5_1/capacitor_5_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C135 charge_pump_reverse_0/capacitors_5_1/capacitor_5_0/buffer_and_gate_0/in1 0 2.57f
C136 charge_pump_reverse_0/nmos_dnw3_0/out2 0 14.9f
C137 charge_pump_reverse_0/capacitors_5_1/capacitor_5_7/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C138 charge_pump_reverse_0/clock_0/clk 0 80f
C139 charge_pump_reverse_0/capacitors_5_1/capacitor_5_7/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C140 charge_pump_reverse_0/capacitors_5_1/capacitor_5_7/buffer_and_gate_0/in1 0 2.57f
C141 charge_pump_reverse_0/capacitors_5_1/capacitor_5_6/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C142 charge_pump_reverse_0/capacitors_5_1/capacitor_5_6/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C143 charge_pump_reverse_0/capacitors_5_1/capacitor_5_6/buffer_and_gate_0/in1 0 2.57f
C144 charge_pump_reverse_0/capacitors_5_1/capacitor_5_5/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C145 charge_pump_reverse_0/capacitors_5_1/capacitor_5_5/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C146 charge_pump_reverse_0/capacitors_5_1/capacitor_5_5/buffer_and_gate_0/in1 0 2.57f
C147 charge_pump_reverse_0/nmos_dnw3_0/clk 0 2.43f
C148 m1_94493_n2143# 0 13.9f
C149 m1_71529_n2069# 0 3.9f
C150 charge_pump_1/clock_0/clk_in 0 13.1f
C151 charge_pump_reverse_0/clock_0/clk_in 0 7.77f
C152 charge_pump_2/nmos_dnw3_0/vs 0 16.4f
C153 charge_pump_2/m1_12174_n760# 0 2.03f
C154 charge_pump_2/clock_0/a_2432_n962# 0 8.68f **FLOATING
C155 charge_pump_2/clock_0/a_2020_n482# 0 2.57f **FLOATING
C156 charge_pump_2/clock_0/a_344_102# 0 2.81f
C157 charge_pump_2/clock_0/a_2402_572# 0 2.17f
C158 charge_pump_2/clock_0/a_344_n986# 0 2.38f
C159 charge_pump_2/clock_0/a_3246_118# 0 6.83f
C160 charge_pump_2/nmos_dnw3_0/vin 0 4.17f
C161 charge_pump_2/nmos_dnw3_0/clkb 0 2.54f
C162 charge_pump_2/capacitors_5_0/capacitor_5_4/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C163 charge_pump_2/capacitors_5_0/capacitor_5_4/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C164 charge_pump_2/capacitors_5_0/capacitor_5_4/buffer_and_gate_0/in1 0 2.57f
C165 charge_pump_2/capacitors_5_0/capacitor_5_3/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C166 charge_pump_2/capacitors_5_0/capacitor_5_3/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C167 charge_pump_2/capacitors_5_0/capacitor_5_3/buffer_and_gate_0/in1 0 2.57f
C168 charge_pump_2/capacitors_5_0/capacitor_5_2/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C169 charge_pump_2/capacitors_5_0/capacitor_5_2/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C170 charge_pump_2/capacitors_5_0/capacitor_5_2/buffer_and_gate_0/in1 0 2.57f
C171 charge_pump_2/capacitors_5_0/capacitor_5_1/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C172 charge_pump_2/capacitors_5_0/capacitor_5_1/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C173 charge_pump_2/capacitors_5_0/capacitor_5_1/buffer_and_gate_0/in1 0 2.57f
C174 m2_91682_21576# 0 5.22f
C175 charge_pump_2/capacitors_5_0/capacitor_5_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C176 charge_pump_2/capacitors_5_0/capacitor_5_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C177 charge_pump_2/capacitors_5_0/capacitor_5_0/buffer_and_gate_0/in1 0 2.57f
C178 charge_pump_2/nmos_dnw3_0/out1 0 15f
C179 charge_pump_2/capacitors_5_0/capacitor_5_7/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C180 charge_pump_2/clock_0/clk 0 78.7f
C181 charge_pump_2/capacitors_5_0/capacitor_5_7/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C182 charge_pump_2/capacitors_5_0/capacitor_5_7/buffer_and_gate_0/in1 0 2.57f
C183 charge_pump_2/capacitors_5_0/capacitor_5_6/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C184 charge_pump_2/capacitors_5_0/capacitor_5_6/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C185 charge_pump_2/capacitors_5_0/capacitor_5_6/buffer_and_gate_0/in1 0 2.57f
C186 charge_pump_2/capacitors_5_0/capacitor_5_5/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C187 charge_pump_2/capacitors_5_0/capacitor_5_5/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C188 charge_pump_2/capacitors_5_0/capacitor_5_5/buffer_and_gate_0/in1 0 2.57f
C189 charge_pump_2/capacitors_5_1/capacitor_5_4/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C190 charge_pump_2/capacitors_5_1/capacitor_5_4/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C191 charge_pump_2/capacitors_5_1/capacitor_5_4/buffer_and_gate_0/in1 0 2.57f
C192 charge_pump_2/capacitors_5_1/capacitor_5_3/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C193 charge_pump_2/capacitors_5_1/capacitor_5_3/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C194 charge_pump_2/capacitors_5_1/capacitor_5_3/buffer_and_gate_0/in1 0 2.57f
C195 charge_pump_2/capacitors_5_1/capacitor_5_2/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C196 charge_pump_2/capacitors_5_1/capacitor_5_2/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C197 charge_pump_2/capacitors_5_1/capacitor_5_2/buffer_and_gate_0/in1 0 2.57f
C198 charge_pump_2/capacitors_5_1/capacitor_5_1/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C199 charge_pump_2/capacitors_5_1/capacitor_5_1/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C200 charge_pump_2/capacitors_5_1/capacitor_5_1/buffer_and_gate_0/in1 0 2.57f
C201 charge_pump_2/capacitors_5_1/capacitor_5_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C202 charge_pump_2/capacitors_5_1/capacitor_5_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C203 charge_pump_2/capacitors_5_1/capacitor_5_0/buffer_and_gate_0/in1 0 2.57f
C204 charge_pump_2/nmos_dnw3_0/out2 0 13.6f
C205 charge_pump_2/capacitors_5_1/capacitor_5_7/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C206 charge_pump_2/clock_0/clkb 0 80.5f
C207 charge_pump_2/capacitors_5_1/capacitor_5_7/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C208 charge_pump_2/capacitors_5_1/capacitor_5_7/buffer_and_gate_0/in1 0 2.57f
C209 charge_pump_2/capacitors_5_1/capacitor_5_6/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C210 charge_pump_2/capacitors_5_1/capacitor_5_6/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C211 charge_pump_2/capacitors_5_1/capacitor_5_6/buffer_and_gate_0/in1 0 2.57f
C212 charge_pump_2/capacitors_5_1/capacitor_5_5/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C213 charge_pump_2/capacitors_5_1/capacitor_5_5/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C214 charge_pump_2/capacitors_5_1/capacitor_5_5/buffer_and_gate_0/in1 0 2.57f
C215 charge_pump_2/nmos_dnw3_0/clk 0 2.76f
C216 charge_pump_1/nmos_dnw3_0/vs 0 16.4f
C217 charge_pump_reverse_1/nmos_dnw3_0/vin 0 3.91f
C218 charge_pump_1/clock_0/a_2432_n962# 0 8.68f **FLOATING
C219 charge_pump_1/clock_0/a_2020_n482# 0 2.57f **FLOATING
C220 charge_pump_1/clock_0/a_344_102# 0 2.81f
C221 charge_pump_1/clock_0/a_2402_572# 0 2.17f
C222 charge_pump_1/clock_0/a_344_n986# 0 2.38f
C223 charge_pump_1/clock_0/a_3246_118# 0 6.83f
C224 charge_pump_1/nmos_dnw3_0/vin 0 4.27f
C225 charge_pump_1/nmos_dnw3_0/clkb 0 2.54f
C226 charge_pump_1/capacitors_5_0/capacitor_5_4/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C227 charge_pump_1/capacitors_5_0/capacitor_5_4/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C228 charge_pump_1/capacitors_5_0/capacitor_5_4/buffer_and_gate_0/in1 0 2.57f
C229 m2_91686_15288# 0 6.65f
C230 charge_pump_1/capacitors_5_0/capacitor_5_3/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C231 charge_pump_1/capacitors_5_0/capacitor_5_3/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C232 charge_pump_1/capacitors_5_0/capacitor_5_3/buffer_and_gate_0/in1 0 2.57f
C233 m2_91690_17386# 0 5.38f
C234 charge_pump_1/capacitors_5_0/capacitor_5_2/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C235 charge_pump_1/capacitors_5_0/capacitor_5_2/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C236 charge_pump_1/capacitors_5_0/capacitor_5_2/buffer_and_gate_0/in1 0 2.57f
C237 charge_pump_1/capacitors_5_0/capacitor_5_1/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C238 charge_pump_1/capacitors_5_0/capacitor_5_1/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C239 charge_pump_1/capacitors_5_0/capacitor_5_1/buffer_and_gate_0/in1 0 2.57f
C240 charge_pump_1/capacitors_5_0/capacitor_5_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C241 charge_pump_1/capacitors_5_0/capacitor_5_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C242 charge_pump_1/capacitors_5_0/capacitor_5_0/buffer_and_gate_0/in1 0 2.57f
C243 charge_pump_1/nmos_dnw3_0/out1 0 15f
C244 charge_pump_1/capacitors_5_0/capacitor_5_7/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C245 charge_pump_1/clock_0/clk 0 78.7f
C246 charge_pump_1/capacitors_5_0/capacitor_5_7/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C247 charge_pump_1/capacitors_5_0/capacitor_5_7/buffer_and_gate_0/in1 0 2.57f
C248 m2_91764_9020# 0 6.43f
C249 charge_pump_1/capacitors_5_0/capacitor_5_6/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C250 charge_pump_1/capacitors_5_0/capacitor_5_6/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C251 charge_pump_1/capacitors_5_0/capacitor_5_6/buffer_and_gate_0/in1 0 2.57f
C252 charge_pump_1/capacitors_5_0/capacitor_5_5/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C253 charge_pump_1/capacitors_5_0/capacitor_5_5/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C254 charge_pump_1/capacitors_5_0/capacitor_5_5/buffer_and_gate_0/in1 0 2.57f
C255 charge_pump_1/capacitors_5_1/capacitor_5_4/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C256 charge_pump_1/capacitors_5_1/capacitor_5_4/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C257 charge_pump_1/capacitors_5_1/capacitor_5_4/buffer_and_gate_0/in1 0 2.57f
C258 charge_pump_1/capacitors_5_1/capacitor_5_3/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C259 charge_pump_1/capacitors_5_1/capacitor_5_3/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C260 charge_pump_1/capacitors_5_1/capacitor_5_3/buffer_and_gate_0/in1 0 2.57f
C261 charge_pump_1/capacitors_5_1/capacitor_5_2/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C262 charge_pump_1/capacitors_5_1/capacitor_5_2/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C263 charge_pump_1/capacitors_5_1/capacitor_5_2/buffer_and_gate_0/in1 0 2.57f
C264 charge_pump_1/capacitors_5_1/capacitor_5_1/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C265 charge_pump_1/capacitors_5_1/capacitor_5_1/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C266 charge_pump_1/capacitors_5_1/capacitor_5_1/buffer_and_gate_0/in1 0 2.57f
C267 charge_pump_1/capacitors_5_1/capacitor_5_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C268 charge_pump_1/capacitors_5_1/capacitor_5_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C269 charge_pump_1/capacitors_5_1/capacitor_5_0/buffer_and_gate_0/in1 0 2.57f
C270 charge_pump_1/nmos_dnw3_0/out2 0 13.6f
C271 charge_pump_1/capacitors_5_1/capacitor_5_7/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C272 charge_pump_1/clock_0/clkb 0 80.5f
C273 charge_pump_1/capacitors_5_1/capacitor_5_7/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C274 charge_pump_1/capacitors_5_1/capacitor_5_7/buffer_and_gate_0/in1 0 2.57f
C275 charge_pump_1/capacitors_5_1/capacitor_5_6/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C276 charge_pump_1/capacitors_5_1/capacitor_5_6/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C277 charge_pump_1/capacitors_5_1/capacitor_5_6/buffer_and_gate_0/in1 0 2.57f
C278 charge_pump_1/capacitors_5_1/capacitor_5_5/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C279 charge_pump_1/capacitors_5_1/capacitor_5_5/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C280 charge_pump_1/capacitors_5_1/capacitor_5_5/buffer_and_gate_0/in1 0 2.57f
C281 charge_pump_1/nmos_dnw3_0/clk 0 2.76f
C282 charge_pump_0/nmos_dnw3_0/vs 0 16.4f
C283 charge_pump_reverse_0/nmos_dnw3_0/vin 0 2.33f
C284 charge_pump_0/clock_0/a_2432_n962# 0 8.68f **FLOATING
C285 charge_pump_0/clock_0/a_2020_n482# 0 2.57f **FLOATING
C286 charge_pump_0/clock_0/a_344_102# 0 2.81f
C287 charge_pump_0/clock_0/a_2402_572# 0 2.17f
C288 charge_pump_0/clock_0/a_344_n986# 0 2.38f
C289 charge_pump_0/clock_0/clk_in 0 15.3f
C290 charge_pump_0/clock_0/a_3246_118# 0 6.83f
C291 charge_pump_0/nmos_dnw3_0/vin 0 2.2f
C292 charge_pump_0/nmos_dnw3_0/clkb 0 2.54f
C293 charge_pump_0/capacitors_5_0/capacitor_5_4/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C294 charge_pump_0/capacitors_5_0/capacitor_5_4/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C295 charge_pump_0/capacitors_5_0/capacitor_5_4/buffer_and_gate_0/in1 0 2.57f
C296 charge_pump_0/capacitors_5_0/capacitor_5_3/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C297 charge_pump_0/capacitors_5_0/capacitor_5_3/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C298 charge_pump_0/capacitors_5_0/capacitor_5_3/buffer_and_gate_0/in1 0 2.57f
C299 charge_pump_0/capacitors_5_0/capacitor_5_2/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C300 charge_pump_0/capacitors_5_0/capacitor_5_2/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C301 charge_pump_0/capacitors_5_0/capacitor_5_2/buffer_and_gate_0/in1 0 2.57f
C302 m2_91690_19482# 0 5.2f
C303 charge_pump_0/capacitors_5_0/capacitor_5_1/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C304 charge_pump_0/capacitors_5_0/capacitor_5_1/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C305 charge_pump_0/capacitors_5_0/capacitor_5_1/buffer_and_gate_0/in1 0 2.57f
C306 charge_pump_0/capacitors_5_0/capacitor_5_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C307 charge_pump_0/capacitors_5_0/capacitor_5_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C308 charge_pump_0/capacitors_5_0/capacitor_5_0/buffer_and_gate_0/in1 0 2.57f
C309 charge_pump_0/nmos_dnw3_0/out1 0 15f
C310 charge_pump_0/capacitors_5_0/capacitor_5_7/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C311 charge_pump_0/clock_0/clk 0 78.7f
C312 charge_pump_0/capacitors_5_0/capacitor_5_7/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C313 VSUBS 0 0.66p
C314 charge_pump_0/capacitors_5_0/capacitor_5_7/buffer_and_gate_0/in1 0 2.57f
C315 charge_pump_0/capacitors_5_0/capacitor_5_6/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C316 charge_pump_0/capacitors_5_0/capacitor_5_6/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C317 charge_pump_0/capacitors_5_0/capacitor_5_6/buffer_and_gate_0/in1 0 2.57f
C318 m2_91760_11118# 0 6.49f
C319 charge_pump_0/capacitors_5_0/capacitor_5_5/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C320 charge_pump_0/capacitors_5_0/capacitor_5_5/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C321 charge_pump_0/capacitors_5_0/capacitor_5_5/buffer_and_gate_0/in1 0 2.57f
C322 m2_91774_13212# 0 6.45f
C323 charge_pump_0/capacitors_5_1/capacitor_5_4/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C324 charge_pump_0/capacitors_5_1/capacitor_5_4/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C325 charge_pump_0/capacitors_5_1/capacitor_5_4/buffer_and_gate_0/in1 0 2.57f
C326 charge_pump_0/capacitors_5_1/capacitor_5_3/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C327 charge_pump_0/capacitors_5_1/capacitor_5_3/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C328 charge_pump_0/capacitors_5_1/capacitor_5_3/buffer_and_gate_0/in1 0 2.57f
C329 charge_pump_0/capacitors_5_1/capacitor_5_2/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C330 charge_pump_0/capacitors_5_1/capacitor_5_2/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C331 charge_pump_0/capacitors_5_1/capacitor_5_2/buffer_and_gate_0/in1 0 2.57f
C332 charge_pump_0/capacitors_5_1/capacitor_5_1/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C333 charge_pump_0/capacitors_5_1/capacitor_5_1/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C334 charge_pump_0/capacitors_5_1/capacitor_5_1/buffer_and_gate_0/in1 0 2.57f
C335 charge_pump_0/capacitors_5_1/capacitor_5_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C336 charge_pump_0/capacitors_5_1/capacitor_5_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C337 charge_pump_0/capacitors_5_1/capacitor_5_0/buffer_and_gate_0/in1 0 2.57f
C338 charge_pump_0/nmos_dnw3_0/out2 0 13.6f
C339 charge_pump_0/capacitors_5_1/capacitor_5_7/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C340 charge_pump_0/clock_0/clkb 0 80.5f
C341 charge_pump_0/capacitors_5_1/capacitor_5_7/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C342 charge_pump_2/clock_0/vdd 0 2.42p
C343 charge_pump_0/capacitors_5_1/capacitor_5_7/buffer_and_gate_0/in1 0 2.57f
C344 charge_pump_0/capacitors_5_1/capacitor_5_6/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C345 charge_pump_0/capacitors_5_1/capacitor_5_6/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C346 charge_pump_0/capacitors_5_1/capacitor_5_6/buffer_and_gate_0/in1 0 2.57f
C347 charge_pump_0/capacitors_5_1/capacitor_5_5/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C348 charge_pump_0/capacitors_5_1/capacitor_5_5/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C349 charge_pump_0/capacitors_5_1/capacitor_5_5/buffer_and_gate_0/in1 0 2.57f
C350 charge_pump_0/nmos_dnw3_0/clk 0 2.76f
.ends

.subckt sky130_fd_pr__nfet_01v8_9LGCGE a_15_n130# a_n561_n130# a_63_n42# a_n989_n42#
+ a_n177_n130# a_n417_n42# a_n465_64# a_255_n42# a_495_64# a_735_n42# a_n129_n42#
+ a_n609_n42# a_111_64# a_447_n42# a_927_n42# a_783_n130# a_n321_n42# a_399_n130#
+ a_n657_64# a_n801_n42# a_687_64# a_n945_n130# a_159_n42# a_639_n42# a_n513_n42#
+ a_n897_n42# a_591_n130# a_n81_64# a_n273_64# a_351_n42# a_207_n130# a_303_64# a_n33_n42#
+ a_831_n42# a_n369_n130# a_n753_n130# a_n849_64# a_n225_n42# a_n705_n42# a_879_64#
+ a_543_n42# VSUBS
X0 a_63_n42# a_15_n130# a_n33_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X1 a_927_n42# a_879_64# a_831_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X2 a_n33_n42# a_n81_64# a_n129_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X3 a_351_n42# a_303_64# a_255_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X4 a_159_n42# a_111_64# a_63_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X5 a_255_n42# a_207_n130# a_159_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X6 a_447_n42# a_399_n130# a_351_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X7 a_543_n42# a_495_64# a_447_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X8 a_735_n42# a_687_64# a_639_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X9 a_831_n42# a_783_n130# a_735_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X10 a_639_n42# a_591_n130# a_543_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X11 a_n321_n42# a_n369_n130# a_n417_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X12 a_n801_n42# a_n849_64# a_n897_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X13 a_n705_n42# a_n753_n130# a_n801_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X14 a_n609_n42# a_n657_64# a_n705_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X15 a_n513_n42# a_n561_n130# a_n609_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X16 a_n417_n42# a_n465_64# a_n513_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X17 a_n225_n42# a_n273_64# a_n321_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X18 a_n129_n42# a_n177_n130# a_n225_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X19 a_n897_n42# a_n945_n130# a_n989_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
.ends

.subckt sky130_fd_pr__pfet_01v8_49FP49 a_63_n42# a_n989_n42# a_n369_n139# a_n753_n139#
+ a_n417_n42# a_687_73# w_n1025_n142# a_255_n42# a_735_n42# a_n81_73# a_n273_73# a_n129_n42#
+ a_15_n139# a_n561_n139# a_303_73# a_n609_n42# a_n177_n139# a_n849_73# a_447_n42#
+ a_927_n42# a_n321_n42# a_879_73# a_n801_n42# a_159_n42# a_639_n42# a_n465_73# a_n513_n42#
+ a_n897_n42# a_783_n139# a_495_73# a_399_n139# a_351_n42# a_n33_n42# a_831_n42# a_n945_n139#
+ a_n225_n42# a_n705_n42# a_111_73# a_591_n139# a_543_n42# a_207_n139# a_n657_73#
+ VSUBS
X0 a_927_n42# a_879_73# a_831_n42# w_n1025_n142# sky130_fd_pr__pfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X1 a_n33_n42# a_n81_73# a_n129_n42# w_n1025_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X2 a_351_n42# a_303_73# a_255_n42# w_n1025_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X3 a_159_n42# a_111_73# a_63_n42# w_n1025_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X4 a_255_n42# a_207_n139# a_159_n42# w_n1025_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X5 a_447_n42# a_399_n139# a_351_n42# w_n1025_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X6 a_543_n42# a_495_73# a_447_n42# w_n1025_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X7 a_639_n42# a_591_n139# a_543_n42# w_n1025_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X8 a_735_n42# a_687_73# a_639_n42# w_n1025_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X9 a_831_n42# a_783_n139# a_735_n42# w_n1025_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X10 a_n801_n42# a_n849_73# a_n897_n42# w_n1025_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X11 a_n513_n42# a_n561_n139# a_n609_n42# w_n1025_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X12 a_n321_n42# a_n369_n139# a_n417_n42# w_n1025_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X13 a_n225_n42# a_n273_73# a_n321_n42# w_n1025_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X14 a_n897_n42# a_n945_n139# a_n989_n42# w_n1025_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.13 ps=1.46 w=0.42 l=0.15
X15 a_n705_n42# a_n753_n139# a_n801_n42# w_n1025_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X16 a_n609_n42# a_n657_73# a_n705_n42# w_n1025_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X17 a_n417_n42# a_n465_73# a_n513_n42# w_n1025_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X18 a_n129_n42# a_n177_n139# a_n225_n42# w_n1025_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X19 a_63_n42# a_15_n139# a_n33_n42# w_n1025_n142# sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
.ends

.subckt capacito7 a_2858_n174# sky130_fd_pr__pfet_01v8_4ZKXAA_0/w_n545_n142# a_5270_n124#
+ m3_7758_166# buffer_and_gate_0/clk sky130_fd_pr__pfet_01v8_49FP49_0/w_n1025_n142#
+ m1_6370_n278# buffer_and_gate_0/gnd buffer_and_gate_0/vdd m1_602_n334# m2_n739_1036#
Xbuffer_digital_0 buffer_and_gate_0/in1 buffer_digital_0/a_116_148# buffer_and_gate_0/vdd
+ buffer_and_gate_0/vdd m2_n739_1036# buffer_and_gate_0/gnd buffer_and_gate_0/gnd
+ buffer_and_gate_0/gnd buffer_digital
Xsky130_fd_pr__pfet_01v8_4ZKXAA_0 m1_6370_n278# m1_6370_n278# buffer_and_gate_0/gnd
+ sky130_fd_pr__pfet_01v8_4ZKXAA_0/w_n545_n142# m1_6370_n278# buffer_and_gate_0/gnd
+ m1_6370_n278# buffer_and_gate_0/gnd m1_6370_n278# buffer_and_gate_0/gnd buffer_and_gate_0/gnd
+ m1_6370_n278# buffer_and_gate_0/gnd m1_6370_n278# m1_6370_n278# buffer_and_gate_0/gnd
+ buffer_and_gate_0/gnd m1_6370_n278# m1_6370_n278# buffer_and_gate_0/gnd m1_6370_n278#
+ buffer_and_gate_0/gnd buffer_and_gate_0/gnd sky130_fd_pr__pfet_01v8_4ZKXAA
Xsky130_fd_pr__nfet_01v8_9LGCGE_0 a_2858_n174# a_2858_n174# buffer_and_gate_0/gnd
+ buffer_and_gate_0/gnd a_2858_n174# buffer_and_gate_0/gnd a_2858_n174# buffer_and_gate_0/gnd
+ a_2858_n174# buffer_and_gate_0/gnd buffer_and_gate_0/gnd buffer_and_gate_0/gnd a_2858_n174#
+ buffer_and_gate_0/gnd buffer_and_gate_0/gnd a_2858_n174# buffer_and_gate_0/gnd a_2858_n174#
+ a_2858_n174# buffer_and_gate_0/gnd a_2858_n174# a_2858_n174# buffer_and_gate_0/gnd
+ buffer_and_gate_0/gnd buffer_and_gate_0/gnd buffer_and_gate_0/gnd a_2858_n174# a_2858_n174#
+ a_2858_n174# buffer_and_gate_0/gnd a_2858_n174# a_2858_n174# buffer_and_gate_0/gnd
+ buffer_and_gate_0/gnd a_2858_n174# a_2858_n174# a_2858_n174# buffer_and_gate_0/gnd
+ buffer_and_gate_0/gnd a_2858_n174# buffer_and_gate_0/gnd buffer_and_gate_0/gnd sky130_fd_pr__nfet_01v8_9LGCGE
Xsky130_fd_pr__pfet_01v8_49FP49_0 m1_602_n334# m1_602_n334# buffer_and_gate_0/gnd
+ buffer_and_gate_0/gnd m1_602_n334# buffer_and_gate_0/gnd sky130_fd_pr__pfet_01v8_49FP49_0/w_n1025_n142#
+ m1_602_n334# m1_602_n334# buffer_and_gate_0/gnd buffer_and_gate_0/gnd m1_602_n334#
+ buffer_and_gate_0/gnd buffer_and_gate_0/gnd buffer_and_gate_0/gnd m1_602_n334# buffer_and_gate_0/gnd
+ buffer_and_gate_0/gnd m1_602_n334# m1_602_n334# m1_602_n334# buffer_and_gate_0/gnd
+ m1_602_n334# m1_602_n334# m1_602_n334# buffer_and_gate_0/gnd m1_602_n334# m1_602_n334#
+ buffer_and_gate_0/gnd buffer_and_gate_0/gnd buffer_and_gate_0/gnd m1_602_n334# m1_602_n334#
+ m1_602_n334# buffer_and_gate_0/gnd m1_602_n334# m1_602_n334# buffer_and_gate_0/gnd
+ buffer_and_gate_0/gnd m1_602_n334# buffer_and_gate_0/gnd buffer_and_gate_0/gnd buffer_and_gate_0/gnd
+ sky130_fd_pr__pfet_01v8_49FP49
Xsky130_fd_pr__nfet_01v8_NJGC45_0 buffer_and_gate_0/gnd a_5270_n124# buffer_and_gate_0/gnd
+ a_5270_n124# a_5270_n124# buffer_and_gate_0/gnd buffer_and_gate_0/gnd a_5270_n124#
+ a_5270_n124# buffer_and_gate_0/gnd a_5270_n124# buffer_and_gate_0/gnd buffer_and_gate_0/gnd
+ buffer_and_gate_0/gnd buffer_and_gate_0/gnd buffer_and_gate_0/gnd a_5270_n124# buffer_and_gate_0/gnd
+ a_5270_n124# a_5270_n124# a_5270_n124# buffer_and_gate_0/gnd sky130_fd_pr__nfet_01v8_NJGC45
Xbuffer_and_gate_0 buffer_and_gate_0/in1 buffer_and_gate_0/clk buffer_and_gate_0/out
+ buffer_and_gate_0/gnd buffer_and_gate_0/vdd buffer_and_gate
X0 buffer_and_gate_0/out m3_7758_166# sky130_fd_pr__cap_mim_m3_1 l=7.99 w=7.97
C0 buffer_and_gate_0/gnd a_2858_n174# 2.03f
C1 buffer_and_gate_0/in1 m2_n739_1036# 2.94f
C2 m3_7758_166# 0 2.32f
C3 buffer_and_gate_0/gnd 0 8.36f
C4 buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C5 buffer_and_gate_0/clk 0 7.7f
C6 buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C7 buffer_and_gate_0/vdd 0 18.2f
C8 a_5270_n124# 0 2.36f
C9 a_2858_n174# 0 4.67f
C10 buffer_and_gate_0/in1 0 2.66f
.ends

.subckt capacitor_8 capacitor_7_0/a_5270_n124# capacitor_7_0/m3_7758_166# capacitor_7_0/buffer_and_gate_0/vdd
+ capacitor_7_0/buffer_and_gate_0/clk capacitor_7_0/a_2858_n174# w_7118_n356# w_1380_n364#
+ VSUBS capacitor_7_0/m2_n739_1036#
Xcapacitor_7_0 capacitor_7_0/a_2858_n174# w_7118_n356# capacitor_7_0/a_5270_n124#
+ capacitor_7_0/m3_7758_166# capacitor_7_0/buffer_and_gate_0/clk w_1380_n364# w_7118_n356#
+ VSUBS capacitor_7_0/buffer_and_gate_0/vdd w_1380_n364# capacitor_7_0/m2_n739_1036#
+ capacito7
C0 capacitor_7_0/m3_7758_166# 0 2.32f
C1 VSUBS 0 8.2f
C2 capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C3 capacitor_7_0/buffer_and_gate_0/clk 0 7.7f
C4 capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C5 capacitor_7_0/buffer_and_gate_0/vdd 0 18.3f
C6 capacitor_7_0/a_5270_n124# 0 2.36f
C7 w_1380_n364# 0 3.28f
C8 capacitor_7_0/a_2858_n174# 0 4.67f
C9 capacitor_7_0/buffer_and_gate_0/in1 0 2.66f
.ends

.subckt capacitors_1 clk1 in1 capacitor_8_0/capacitor_7_0/a_2858_n174# capacitor_8_0/capacitor_7_0/a_5270_n124#
+ capacitor_8_0/capacitor_7_0/buffer_and_gate_0/clk capacitor_8_0/capacitor_7_0/buffer_and_gate_0/vdd
+ m1_7096_n308# capacitor_8_0/w_1380_n364# VSUBS
Xcapacitor_8_0 capacitor_8_0/capacitor_7_0/a_5270_n124# clk1 capacitor_8_0/capacitor_7_0/buffer_and_gate_0/vdd
+ capacitor_8_0/capacitor_7_0/buffer_and_gate_0/clk capacitor_8_0/capacitor_7_0/a_2858_n174#
+ m1_7096_n308# capacitor_8_0/w_1380_n364# VSUBS in1 capacitor_8
C0 VSUBS capacitor_8_0/capacitor_7_0/buffer_and_gate_0/vdd 2.83f
C1 clk1 0 2.38f
C2 VSUBS 0 8.2f
C3 capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C4 capacitor_8_0/capacitor_7_0/buffer_and_gate_0/clk 0 8.5f
C5 capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C6 capacitor_8_0/capacitor_7_0/buffer_and_gate_0/vdd 0 18.3f
C7 capacitor_8_0/capacitor_7_0/a_5270_n124# 0 2.36f
C8 capacitor_8_0/w_1380_n364# 0 3.28f
C9 capacitor_8_0/capacitor_7_0/a_2858_n174# 0 4.67f
C10 capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 0 2.66f
.ends

.subckt sky130_fd_pr__pfet_01v8_E9H44Q a_15_n42# a_n15_n68# w_n109_n104# a_n73_n42#
+ VSUBS
X0 a_15_n42# a_n15_n68# a_n73_n42# w_n109_n104# sky130_fd_pr__pfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
.ends

.subckt sky130_fd_pr__pfet_01v8_9AYYDL a_n158_n300# w_n194_n362# a_100_n300# a_n100_n326#
+ VSUBS
X0 a_100_n300# a_n100_n326# a_n158_n300# w_n194_n362# sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.87 ps=6.58 w=3 l=1
.ends

.subckt pmos_cp1 a_168_22# m1_532_58# w_n14_n142# a_424_18# m1_14_56# VSUBS
Xsky130_fd_pr__pfet_01v8_E9H44Q_0 w_n14_n142# a_168_22# w_n14_n142# a_424_18# VSUBS
+ sky130_fd_pr__pfet_01v8_E9H44Q
Xsky130_fd_pr__pfet_01v8_E9H44Q_1 a_168_22# a_424_18# w_n14_n142# w_n14_n142# VSUBS
+ sky130_fd_pr__pfet_01v8_E9H44Q
Xsky130_fd_pr__pfet_01v8_9AYYDL_0 m1_14_56# w_n14_n142# w_n14_n142# a_168_22# VSUBS
+ sky130_fd_pr__pfet_01v8_9AYYDL
Xsky130_fd_pr__pfet_01v8_9AYYDL_1 w_n14_n142# w_n14_n142# m1_532_58# a_424_18# VSUBS
+ sky130_fd_pr__pfet_01v8_9AYYDL
C0 w_n14_n142# VSUBS 2.47f
.ends

.subckt charge_pump1 clk_in input1 input2 vdd in5 in6 in8 m1_12464_n576# a_3340_18086#
+ in3 in4 gnd nmos_dnw3_0/vs in1 in2 in7
Xsky130_fd_pr__cap_mim_m3_1_MH6KF8_4 nmos_dnw3_0/clk clock_0/clk gnd sky130_fd_pr__cap_mim_m3_1_MH6KF8
Xsky130_fd_pr__cap_mim_m3_1_MH6KF8_5 nmos_dnw3_0/clkb clock_0/clkb gnd sky130_fd_pr__cap_mim_m3_1_MH6KF8
Xnmos_dnw3_0 nmos_dnw3_0/vs input1 input2 nmos_dnw3_0/clk nmos_dnw3_0/clkb nmos_dnw3_0/vs
+ gnd nmos_dnw3
Xclock_0 clk_in vdd gnd clock_0/clk clock_0/clkb clock
Xcapacitor_8_0 vdd input1 vdd clock_0/clk vdd vdd vdd gnd in8 capacitor_8
Xcapacitor_8_1 vdd input2 vdd clock_0/clkb vdd vdd vdd gnd in8 capacitor_8
Xcapacitors_1_0 input1 in1 vdd vdd clock_0/clk vdd vdd vdd gnd capacitors_1
Xcapacitors_1_1 input2 in1 vdd vdd clock_0/clkb vdd vdd vdd gnd capacitors_1
Xcapacitors_1_2 input1 in2 vdd vdd clock_0/clk vdd vdd vdd gnd capacitors_1
Xsky130_fd_pr__pfet_01v8_4RPJ49_0 gnd vdd vdd gnd gnd vdd vdd vdd gnd vdd gnd gnd
+ vdd gnd gnd gnd vdd vdd vdd vdd gnd vdd gnd gnd gnd gnd gnd gnd gnd vdd gnd vdd
+ gnd gnd vdd gnd gnd vdd vdd gnd vdd gnd gnd vdd gnd gnd vdd vdd gnd gnd vdd vdd
+ vdd gnd gnd vdd vdd gnd gnd vdd vdd gnd vdd gnd vdd gnd gnd gnd vdd gnd gnd gnd
+ vdd vdd gnd gnd vdd vdd gnd gnd vdd vdd gnd gnd gnd vdd vdd vdd vdd vdd vdd vdd
+ vdd vdd gnd gnd vdd vdd vdd gnd vdd vdd vdd vdd vdd gnd vdd vdd gnd vdd vdd gnd
+ gnd gnd gnd gnd vdd vdd vdd gnd vdd vdd gnd vdd gnd vdd vdd vdd gnd gnd vdd vdd
+ gnd vdd vdd vdd vdd gnd vdd gnd gnd gnd vdd vdd vdd gnd gnd gnd gnd vdd gnd gnd
+ gnd vdd gnd gnd gnd gnd vdd gnd gnd vdd vdd sky130_fd_pr__pfet_01v8_4RPJ49
Xcapacitors_1_3 input1 in3 vdd vdd clock_0/clk vdd vdd vdd gnd capacitors_1
Xsky130_fd_pr__pfet_01v8_4RPJ49_1 gnd vdd vdd gnd gnd vdd vdd vdd gnd vdd gnd gnd
+ vdd gnd gnd gnd vdd vdd vdd vdd gnd vdd gnd gnd gnd gnd gnd gnd gnd vdd gnd vdd
+ gnd gnd vdd gnd gnd vdd vdd gnd vdd gnd gnd vdd gnd gnd vdd vdd gnd gnd vdd vdd
+ vdd gnd gnd vdd vdd gnd gnd vdd vdd gnd vdd gnd vdd gnd gnd gnd vdd gnd gnd gnd
+ vdd vdd gnd gnd vdd vdd gnd gnd vdd vdd gnd gnd gnd vdd vdd vdd vdd vdd vdd vdd
+ vdd vdd gnd gnd vdd vdd vdd gnd vdd vdd vdd vdd vdd gnd vdd vdd gnd vdd vdd gnd
+ gnd gnd gnd gnd vdd vdd vdd gnd vdd vdd gnd vdd gnd vdd vdd vdd gnd gnd vdd vdd
+ gnd vdd vdd vdd vdd gnd vdd gnd gnd gnd vdd vdd vdd gnd gnd gnd gnd vdd gnd gnd
+ gnd vdd gnd gnd gnd gnd vdd gnd gnd vdd vdd sky130_fd_pr__pfet_01v8_4RPJ49
Xcapacitors_1_4 input2 in2 vdd vdd clock_0/clkb vdd vdd vdd gnd capacitors_1
Xcapacitors_1_5 input2 in3 vdd vdd clock_0/clkb vdd vdd vdd gnd capacitors_1
Xcapacitors_1_6 input1 in4 vdd vdd clock_0/clk vdd vdd vdd gnd capacitors_1
Xcapacitors_1_7 input1 in5 vdd vdd clock_0/clk vdd vdd vdd gnd capacitors_1
Xcapacitors_1_8 input1 in6 vdd vdd clock_0/clk vdd vdd vdd gnd capacitors_1
Xcapacitors_1_9 input1 in7 vdd vdd clock_0/clk vdd vdd vdd gnd capacitors_1
Xpmos_cp1_0 m1_12659_300# input2 m1_12464_n576# m1_4341_n519# input1 gnd pmos_cp1
Xsky130_fd_pr__nfet_01v8_NJGC8F_0 vdd gnd gnd vdd vdd gnd gnd vdd gnd vdd gnd gnd
+ vdd gnd gnd gnd vdd gnd vdd vdd gnd vdd vdd vdd vdd gnd vdd vdd gnd vdd vdd gnd
+ gnd gnd gnd gnd vdd gnd gnd vdd gnd gnd gnd vdd gnd gnd vdd gnd gnd gnd vdd vdd
+ gnd gnd vdd gnd gnd vdd gnd gnd gnd vdd vdd vdd gnd gnd gnd gnd vdd gnd vdd gnd
+ vdd gnd gnd vdd gnd vdd vdd vdd vdd vdd vdd gnd gnd gnd gnd gnd vdd gnd gnd vdd
+ vdd gnd vdd vdd vdd vdd gnd vdd gnd gnd gnd gnd gnd vdd vdd vdd vdd gnd vdd vdd
+ vdd vdd gnd vdd gnd vdd vdd gnd gnd vdd gnd gnd vdd vdd vdd gnd gnd vdd gnd gnd
+ gnd vdd vdd gnd vdd vdd vdd gnd vdd vdd gnd gnd gnd vdd vdd vdd gnd vdd vdd vdd
+ vdd vdd vdd gnd vdd gnd vdd gnd gnd gnd sky130_fd_pr__nfet_01v8_NJGC8F
Xcapacitors_1_10 input2 in7 vdd vdd clock_0/clkb vdd vdd vdd gnd capacitors_1
Xcapacitors_1_11 input2 in6 vdd vdd clock_0/clkb vdd vdd vdd gnd capacitors_1
Xsky130_fd_pr__nfet_01v8_NJGC8F_1 vdd gnd gnd vdd vdd gnd gnd vdd gnd vdd gnd gnd
+ vdd gnd gnd gnd vdd gnd vdd vdd gnd vdd vdd vdd vdd gnd vdd vdd gnd vdd vdd gnd
+ gnd gnd gnd gnd vdd gnd gnd vdd gnd gnd gnd vdd gnd gnd vdd gnd gnd gnd vdd vdd
+ gnd gnd vdd gnd gnd vdd gnd gnd gnd vdd vdd vdd gnd gnd gnd gnd vdd gnd vdd gnd
+ vdd gnd gnd vdd gnd vdd vdd vdd vdd vdd vdd gnd gnd gnd gnd gnd vdd gnd gnd vdd
+ vdd gnd vdd vdd vdd vdd gnd vdd gnd gnd gnd gnd gnd vdd vdd vdd vdd gnd vdd vdd
+ vdd vdd gnd vdd gnd vdd vdd gnd gnd vdd gnd gnd vdd vdd vdd gnd gnd vdd gnd gnd
+ gnd vdd vdd gnd vdd vdd vdd gnd vdd vdd gnd gnd gnd vdd vdd vdd gnd vdd vdd vdd
+ vdd vdd vdd gnd vdd gnd vdd gnd gnd gnd sky130_fd_pr__nfet_01v8_NJGC8F
Xcapacitors_1_13 input2 in4 vdd vdd clock_0/clkb vdd vdd vdd gnd capacitors_1
Xcapacitors_1_12 input2 in5 vdd vdd clock_0/clkb vdd vdd vdd gnd capacitors_1
Xsky130_fd_pr__cap_mim_m3_1_MH6KF8_0 clock_0/clkb input2 gnd sky130_fd_pr__cap_mim_m3_1_MH6KF8
Xsky130_fd_pr__cap_mim_m3_1_MH6KF8_1 clock_0/clk input1 gnd sky130_fd_pr__cap_mim_m3_1_MH6KF8
Xsky130_fd_pr__cap_mim_m3_1_MH6KF8_3 m1_12659_300# clock_0/clkb gnd sky130_fd_pr__cap_mim_m3_1_MH6KF8
Xsky130_fd_pr__cap_mim_m3_1_MH6KF8_2 m1_4341_n519# clock_0/clk gnd sky130_fd_pr__cap_mim_m3_1_MH6KF8
C0 gnd clock_0/clk 2.49f
C1 vdd clock_0/clkb 26f
C2 m1_12464_n576# clock_0/clk 2.31f
C3 gnd input1 8.5f
C4 vdd clock_0/clk 32f
C5 vdd gnd 0.171p
C6 clock_0/clk nmos_dnw3_0/vs 2.19f
C7 gnd input2 8.88f
C8 vdd input1 26.8f
C9 input1 input2 3.06f
C10 vdd input2 26.5f
C11 vdd nmos_dnw3_0/vs 9.13f
C12 m1_12464_n576# clock_0/clkb 2.21f
C13 input1 0 22.5f
C14 input2 0 22.2f
C15 capacitors_1_12/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C16 capacitors_1_12/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C17 capacitors_1_12/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 0 2.66f
C18 capacitors_1_13/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C19 capacitors_1_13/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C20 capacitors_1_13/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 0 2.66f
C21 capacitors_1_11/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C22 capacitors_1_11/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C23 capacitors_1_11/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 0 2.66f
C24 capacitors_1_10/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C25 capacitors_1_10/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C26 capacitors_1_10/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 0 2.66f
C27 m1_4341_n519# 0 3.77f
C28 m1_12659_300# 0 2.54f
C29 m1_12464_n576# 0 4.25f
C30 capacitors_1_9/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C31 capacitors_1_9/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C32 capacitors_1_9/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 0 2.66f
C33 capacitors_1_8/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C34 capacitors_1_8/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C35 capacitors_1_8/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 0 2.66f
C36 capacitors_1_7/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C37 capacitors_1_7/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C38 capacitors_1_7/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 0 2.66f
C39 capacitors_1_6/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C40 capacitors_1_6/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C41 capacitors_1_6/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 0 2.66f
C42 capacitors_1_5/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C43 capacitors_1_5/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C44 capacitors_1_5/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 0 2.66f
C45 capacitors_1_4/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C46 capacitors_1_4/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C47 capacitors_1_4/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 0 2.66f
C48 capacitors_1_3/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C49 capacitors_1_3/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C50 capacitors_1_3/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 0 2.66f
C51 capacitors_1_2/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C52 capacitors_1_2/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C53 capacitors_1_2/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 0 2.66f
C54 capacitors_1_1/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C55 capacitors_1_1/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C56 capacitors_1_1/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 0 2.66f
C57 capacitors_1_0/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C58 capacitors_1_0/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C59 capacitors_1_0/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 0 2.66f
C60 capacitor_8_1/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C61 clock_0/clkb 0 86.1f
C62 capacitor_8_1/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C63 capacitor_8_1/capacitor_7_0/buffer_and_gate_0/in1 0 2.66f
C64 gnd 0 48.9f
C65 capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C66 clock_0/clk 0 85.5f
C67 capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C68 vdd 0 0.458p
C69 capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 0 2.66f
C70 clock_0/a_2432_n962# 0 8.68f **FLOATING
C71 clock_0/a_2020_n482# 0 2.57f **FLOATING
C72 clock_0/a_344_102# 0 2.81f
C73 clock_0/a_2402_572# 0 2.17f
C74 clock_0/a_344_n986# 0 2.38f
C75 clock_0/a_3246_118# 0 6.83f
C76 nmos_dnw3_0/clkb 0 2.34f
C77 nmos_dnw3_0/vs 0 10.4f
.ends

.subckt charge_pump1_reverse input1 input2 in1 in5 in6 in8 vdd m1_12464_n576# clock_1/clk_in
+ a_3340_18086# gnd in4 in3 nmos_dnw3_0/vs in7 in2
Xsky130_fd_pr__cap_mim_m3_1_MH6KF8_4 nmos_dnw3_0/clk clock_1/clkb gnd sky130_fd_pr__cap_mim_m3_1_MH6KF8
Xsky130_fd_pr__cap_mim_m3_1_MH6KF8_5 nmos_dnw3_0/clkb clock_1/clk gnd sky130_fd_pr__cap_mim_m3_1_MH6KF8
Xnmos_dnw3_0 nmos_dnw3_0/vs input1 input2 nmos_dnw3_0/clk nmos_dnw3_0/clkb nmos_dnw3_0/vs
+ gnd nmos_dnw3
Xclock_1 clock_1/clk_in vdd gnd clock_1/clk clock_1/clkb clock
Xcapacitor_8_0 vdd input1 vdd clock_1/clkb vdd vdd vdd gnd in8 capacitor_8
Xcapacitor_8_1 vdd input2 vdd clock_1/clk vdd vdd vdd gnd in8 capacitor_8
Xcapacitors_1_0 input1 in1 vdd vdd clock_1/clkb vdd vdd vdd gnd capacitors_1
Xcapacitors_1_1 input2 in1 vdd vdd clock_1/clk vdd vdd vdd gnd capacitors_1
Xcapacitors_1_2 input1 in2 vdd vdd clock_1/clkb vdd vdd vdd gnd capacitors_1
Xsky130_fd_pr__pfet_01v8_4RPJ49_0 gnd vdd vdd gnd gnd vdd vdd vdd gnd vdd gnd gnd
+ vdd gnd gnd gnd vdd vdd vdd vdd gnd vdd gnd gnd gnd gnd gnd gnd gnd vdd gnd vdd
+ gnd gnd vdd gnd gnd vdd vdd gnd vdd gnd gnd vdd gnd gnd vdd vdd gnd gnd vdd vdd
+ vdd gnd gnd vdd vdd gnd gnd vdd vdd gnd vdd gnd vdd gnd gnd gnd vdd gnd gnd gnd
+ vdd vdd gnd gnd vdd vdd gnd gnd vdd vdd gnd gnd gnd vdd vdd vdd vdd vdd vdd vdd
+ vdd vdd gnd gnd vdd vdd vdd gnd vdd vdd vdd vdd vdd gnd vdd vdd gnd vdd vdd gnd
+ gnd gnd gnd gnd vdd vdd vdd gnd vdd vdd gnd vdd gnd vdd vdd vdd gnd gnd vdd vdd
+ gnd vdd vdd vdd vdd gnd vdd gnd gnd gnd vdd vdd vdd gnd gnd gnd gnd vdd gnd gnd
+ gnd vdd gnd gnd gnd gnd vdd gnd gnd vdd vdd sky130_fd_pr__pfet_01v8_4RPJ49
Xsky130_fd_pr__pfet_01v8_4RPJ49_1 gnd vdd vdd gnd gnd vdd vdd vdd gnd vdd gnd gnd
+ vdd gnd gnd gnd vdd vdd vdd vdd gnd vdd gnd gnd gnd gnd gnd gnd gnd vdd gnd vdd
+ gnd gnd vdd gnd gnd vdd vdd gnd vdd gnd gnd vdd gnd gnd vdd vdd gnd gnd vdd vdd
+ vdd gnd gnd vdd vdd gnd gnd vdd vdd gnd vdd gnd vdd gnd gnd gnd vdd gnd gnd gnd
+ vdd vdd gnd gnd vdd vdd gnd gnd vdd vdd gnd gnd gnd vdd vdd vdd vdd vdd vdd vdd
+ vdd vdd gnd gnd vdd vdd vdd gnd vdd vdd vdd vdd vdd gnd vdd vdd gnd vdd vdd gnd
+ gnd gnd gnd gnd vdd vdd vdd gnd vdd vdd gnd vdd gnd vdd vdd vdd gnd gnd vdd vdd
+ gnd vdd vdd vdd vdd gnd vdd gnd gnd gnd vdd vdd vdd gnd gnd gnd gnd vdd gnd gnd
+ gnd vdd gnd gnd gnd gnd vdd gnd gnd vdd vdd sky130_fd_pr__pfet_01v8_4RPJ49
Xcapacitors_1_3 input1 in3 vdd vdd clock_1/clkb vdd vdd vdd gnd capacitors_1
Xcapacitors_1_4 input2 in2 vdd vdd clock_1/clk vdd vdd vdd gnd capacitors_1
Xcapacitors_1_5 input2 in3 vdd vdd clock_1/clk vdd vdd vdd gnd capacitors_1
Xcapacitors_1_6 input1 in4 vdd vdd clock_1/clkb vdd vdd vdd gnd capacitors_1
Xcapacitors_1_7 input1 in5 vdd vdd clock_1/clkb vdd vdd vdd gnd capacitors_1
Xcapacitors_1_8 input1 in6 vdd vdd clock_1/clkb vdd vdd vdd gnd capacitors_1
Xcapacitors_1_9 input1 in7 vdd vdd clock_1/clkb vdd vdd vdd gnd capacitors_1
Xpmos_cp1_0 m1_12659_300# input2 m1_12464_n576# m1_4341_n519# input1 gnd pmos_cp1
Xsky130_fd_pr__nfet_01v8_NJGC8F_0 vdd gnd gnd vdd vdd gnd gnd vdd gnd vdd gnd gnd
+ vdd gnd gnd gnd vdd gnd vdd vdd gnd vdd vdd vdd vdd gnd vdd vdd gnd vdd vdd gnd
+ gnd gnd gnd gnd vdd gnd gnd vdd gnd gnd gnd vdd gnd gnd vdd gnd gnd gnd vdd vdd
+ gnd gnd vdd gnd gnd vdd gnd gnd gnd vdd vdd vdd gnd gnd gnd gnd vdd gnd vdd gnd
+ vdd gnd gnd vdd gnd vdd vdd vdd vdd vdd vdd gnd gnd gnd gnd gnd vdd gnd gnd vdd
+ vdd gnd vdd vdd vdd vdd gnd vdd gnd gnd gnd gnd gnd vdd vdd vdd vdd gnd vdd vdd
+ vdd vdd gnd vdd gnd vdd vdd gnd gnd vdd gnd gnd vdd vdd vdd gnd gnd vdd gnd gnd
+ gnd vdd vdd gnd vdd vdd vdd gnd vdd vdd gnd gnd gnd vdd vdd vdd gnd vdd vdd vdd
+ vdd vdd vdd gnd vdd gnd vdd gnd gnd gnd sky130_fd_pr__nfet_01v8_NJGC8F
Xcapacitors_1_10 input2 in7 vdd vdd clock_1/clk vdd vdd vdd gnd capacitors_1
Xcapacitors_1_11 input2 in6 vdd vdd clock_1/clk vdd vdd vdd gnd capacitors_1
Xsky130_fd_pr__nfet_01v8_NJGC8F_1 vdd gnd gnd vdd vdd gnd gnd vdd gnd vdd gnd gnd
+ vdd gnd gnd gnd vdd gnd vdd vdd gnd vdd vdd vdd vdd gnd vdd vdd gnd vdd vdd gnd
+ gnd gnd gnd gnd vdd gnd gnd vdd gnd gnd gnd vdd gnd gnd vdd gnd gnd gnd vdd vdd
+ gnd gnd vdd gnd gnd vdd gnd gnd gnd vdd vdd vdd gnd gnd gnd gnd vdd gnd vdd gnd
+ vdd gnd gnd vdd gnd vdd vdd vdd vdd vdd vdd gnd gnd gnd gnd gnd vdd gnd gnd vdd
+ vdd gnd vdd vdd vdd vdd gnd vdd gnd gnd gnd gnd gnd vdd vdd vdd vdd gnd vdd vdd
+ vdd vdd gnd vdd gnd vdd vdd gnd gnd vdd gnd gnd vdd vdd vdd gnd gnd vdd gnd gnd
+ gnd vdd vdd gnd vdd vdd vdd gnd vdd vdd gnd gnd gnd vdd vdd vdd gnd vdd vdd vdd
+ vdd vdd vdd gnd vdd gnd vdd gnd gnd gnd sky130_fd_pr__nfet_01v8_NJGC8F
Xcapacitors_1_13 input2 in4 vdd vdd clock_1/clk vdd vdd vdd gnd capacitors_1
Xcapacitors_1_12 input2 in5 vdd vdd clock_1/clk vdd vdd vdd gnd capacitors_1
Xsky130_fd_pr__cap_mim_m3_1_MH6KF8_0 clock_1/clk input2 gnd sky130_fd_pr__cap_mim_m3_1_MH6KF8
Xsky130_fd_pr__cap_mim_m3_1_MH6KF8_1 clock_1/clkb input1 gnd sky130_fd_pr__cap_mim_m3_1_MH6KF8
Xsky130_fd_pr__cap_mim_m3_1_MH6KF8_3 m1_12659_300# clock_1/clk gnd sky130_fd_pr__cap_mim_m3_1_MH6KF8
Xsky130_fd_pr__cap_mim_m3_1_MH6KF8_2 m1_4341_n519# clock_1/clkb gnd sky130_fd_pr__cap_mim_m3_1_MH6KF8
C0 nmos_dnw3_0/vs clock_1/clkb 2.22f
C1 nmos_dnw3_0/vs vdd 9.23f
C2 input2 vdd 26.5f
C3 input1 input2 3.06f
C4 clock_1/clkb vdd 31.8f
C5 m1_12464_n576# clock_1/clkb 2.02f
C6 gnd input2 8.27f
C7 input1 vdd 26.5f
C8 gnd clock_1/clkb 2.85f
C9 gnd vdd 0.166p
C10 input1 gnd 8.5f
C11 clock_1/clk vdd 28.4f
C12 input1 0 22.9f
C13 input2 0 22.4f
C14 capacitors_1_12/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C15 capacitors_1_12/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C16 capacitors_1_12/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 0 2.66f
C17 capacitors_1_13/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C18 capacitors_1_13/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C19 capacitors_1_13/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 0 2.66f
C20 capacitors_1_11/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C21 capacitors_1_11/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C22 capacitors_1_11/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 0 2.66f
C23 capacitors_1_10/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C24 capacitors_1_10/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C25 capacitors_1_10/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 0 2.66f
C26 m1_4341_n519# 0 3.86f
C27 m1_12659_300# 0 2.73f
C28 m1_12464_n576# 0 4.64f
C29 capacitors_1_9/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C30 capacitors_1_9/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C31 capacitors_1_9/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 0 2.66f
C32 capacitors_1_8/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C33 capacitors_1_8/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C34 capacitors_1_8/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 0 2.66f
C35 capacitors_1_7/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C36 capacitors_1_7/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C37 capacitors_1_7/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 0 2.66f
C38 capacitors_1_6/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C39 capacitors_1_6/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C40 capacitors_1_6/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 0 2.66f
C41 capacitors_1_5/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C42 capacitors_1_5/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C43 capacitors_1_5/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 0 2.66f
C44 capacitors_1_4/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C45 capacitors_1_4/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C46 capacitors_1_4/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 0 2.66f
C47 capacitors_1_3/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C48 capacitors_1_3/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C49 capacitors_1_3/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 0 2.66f
C50 capacitors_1_2/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C51 capacitors_1_2/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C52 capacitors_1_2/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 0 2.66f
C53 capacitors_1_1/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C54 capacitors_1_1/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C55 capacitors_1_1/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 0 2.66f
C56 capacitors_1_0/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C57 capacitors_1_0/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C58 capacitors_1_0/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 0 2.66f
C59 capacitor_8_1/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C60 clock_1/clk 0 88.1f
C61 capacitor_8_1/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C62 capacitor_8_1/capacitor_7_0/buffer_and_gate_0/in1 0 2.66f
C63 gnd 0 54.5f
C64 capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C65 clock_1/clkb 0 96.8f
C66 capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C67 vdd 0 0.462p
C68 capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 0 2.66f
C69 clock_1/a_2432_n962# 0 8.68f **FLOATING
C70 clock_1/a_2020_n482# 0 2.57f **FLOATING
C71 clock_1/a_344_102# 0 2.81f
C72 clock_1/a_2402_572# 0 2.17f
C73 clock_1/a_344_n986# 0 2.38f
C74 clock_1/a_3246_118# 0 6.83f
C75 nmos_dnw3_0/clkb 0 2.01f
C76 nmos_dnw3_0/vs 0 10.4f
.ends

.subckt CP1_5_stage charge_pump1_2/vdd charge_pump1_2/in8 charge_pump1_2/in1 charge_pump1_2/in2
+ charge_pump1_2/m1_12464_n576# charge_pump1_2/in3 charge_pump1_reverse_0/nmos_dnw3_0/vs
+ charge_pump1_2/in4 charge_pump1_1/nmos_dnw3_0/vs charge_pump1_0/clk_in charge_pump1_2/in5
+ charge_pump1_2/in6 charge_pump1_0/nmos_dnw3_0/vs charge_pump1_2/in7 charge_pump1_reverse_1/nmos_dnw3_0/vs
+ charge_pump1_2/nmos_dnw3_0/vs VSUBS
Xcharge_pump1_0 charge_pump1_0/clk_in charge_pump1_0/input1 charge_pump1_0/input2
+ charge_pump1_2/vdd charge_pump1_2/in5 charge_pump1_2/in6 charge_pump1_2/in8 charge_pump1_reverse_0/nmos_dnw3_0/vs
+ VSUBS charge_pump1_2/in3 charge_pump1_2/in4 VSUBS charge_pump1_0/nmos_dnw3_0/vs
+ charge_pump1_2/in1 charge_pump1_2/in2 charge_pump1_2/in7 charge_pump1
Xcharge_pump1_1 charge_pump1_1/clk_in charge_pump1_1/input1 charge_pump1_1/input2
+ charge_pump1_2/vdd charge_pump1_2/in5 charge_pump1_2/in6 charge_pump1_2/in8 charge_pump1_reverse_1/nmos_dnw3_0/vs
+ charge_pump1_1/a_3340_18086# charge_pump1_2/in3 charge_pump1_2/in4 VSUBS charge_pump1_1/nmos_dnw3_0/vs
+ charge_pump1_2/in1 charge_pump1_2/in2 charge_pump1_2/in7 charge_pump1
Xcharge_pump1_2 charge_pump1_2/clk_in charge_pump1_2/input1 charge_pump1_2/input2
+ charge_pump1_2/vdd charge_pump1_2/in5 charge_pump1_2/in6 charge_pump1_2/in8 charge_pump1_2/m1_12464_n576#
+ charge_pump1_2/a_3340_18086# charge_pump1_2/in3 charge_pump1_2/in4 VSUBS charge_pump1_2/nmos_dnw3_0/vs
+ charge_pump1_2/in1 charge_pump1_2/in2 charge_pump1_2/in7 charge_pump1
Xbuffer_digital_0 m1_24170_n2398# buffer_digital_0/a_116_148# charge_pump1_2/vdd charge_pump1_2/vdd
+ charge_pump1_0/clk_in VSUBS VSUBS VSUBS buffer_digital
Xcharge_pump1_reverse_0 charge_pump1_reverse_0/input1 charge_pump1_reverse_0/input2
+ charge_pump1_2/in8 charge_pump1_2/in4 charge_pump1_2/in3 charge_pump1_2/in1 charge_pump1_2/vdd
+ charge_pump1_1/nmos_dnw3_0/vs charge_pump1_reverse_0/clock_1/clk_in VSUBS VSUBS
+ charge_pump1_2/in5 charge_pump1_2/in6 charge_pump1_reverse_0/nmos_dnw3_0/vs charge_pump1_2/in2
+ charge_pump1_2/in7 charge_pump1_reverse
Xbuffer_digital_1 charge_pump1_reverse_0/clock_1/clk_in m1_24170_n2398# charge_pump1_2/vdd
+ charge_pump1_2/vdd m1_24170_n2398# VSUBS VSUBS VSUBS buffer_digital
Xcharge_pump1_reverse_1 charge_pump1_reverse_1/input1 charge_pump1_reverse_1/input2
+ charge_pump1_2/in8 charge_pump1_2/in4 charge_pump1_2/in3 charge_pump1_2/in1 charge_pump1_2/vdd
+ charge_pump1_2/nmos_dnw3_0/vs charge_pump1_reverse_1/clock_1/clk_in VSUBS VSUBS
+ charge_pump1_2/in5 charge_pump1_2/in6 charge_pump1_reverse_1/nmos_dnw3_0/vs charge_pump1_2/in2
+ charge_pump1_2/in7 charge_pump1_reverse
X0 a_73934_n2624# charge_pump1_1/clk_in charge_pump1_2/vdd charge_pump1_2/vdd sky130_fd_pr__pfet_01v8 ad=0.365 pd=3.1 as=0.365 ps=3.1 w=1.26 l=0.15
X1 a_100152_n2424# a_99934_n2424# charge_pump1_2/vdd charge_pump1_2/vdd sky130_fd_pr__pfet_01v8 ad=0.365 pd=3.1 as=0.365 ps=3.1 w=1.26 l=0.15
X2 charge_pump1_reverse_1/clock_1/clk_in a_80522_n2634# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X3 charge_pump1_reverse_1/clock_1/clk_in a_80522_n2634# charge_pump1_2/vdd charge_pump1_2/vdd sky130_fd_pr__pfet_01v8 ad=0.365 pd=3.1 as=0.365 ps=3.1 w=1.26 l=0.15
X4 a_48152_n2524# a_47934_n2524# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X5 a_54522_n2534# a_48152_n2524# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X6 a_48152_n2524# a_47934_n2524# charge_pump1_2/vdd charge_pump1_2/vdd sky130_fd_pr__pfet_01v8 ad=0.365 pd=3.1 as=0.365 ps=3.1 w=1.26 l=0.15
X7 a_54522_n2534# a_48152_n2524# charge_pump1_2/vdd charge_pump1_2/vdd sky130_fd_pr__pfet_01v8 ad=0.365 pd=3.1 as=0.365 ps=3.1 w=1.26 l=0.15
X8 a_106522_n2434# a_100152_n2424# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X9 a_47934_n2524# charge_pump1_reverse_0/clock_1/clk_in VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X10 a_106522_n2434# a_100152_n2424# charge_pump1_2/vdd charge_pump1_2/vdd sky130_fd_pr__pfet_01v8 ad=0.365 pd=3.1 as=0.365 ps=3.1 w=1.26 l=0.15
X11 a_47934_n2524# charge_pump1_reverse_0/clock_1/clk_in charge_pump1_2/vdd charge_pump1_2/vdd sky130_fd_pr__pfet_01v8 ad=0.365 pd=3.1 as=0.365 ps=3.1 w=1.26 l=0.15
X12 charge_pump1_1/clk_in a_54522_n2534# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X13 charge_pump1_1/clk_in a_54522_n2534# charge_pump1_2/vdd charge_pump1_2/vdd sky130_fd_pr__pfet_01v8 ad=0.365 pd=3.1 as=0.365 ps=3.1 w=1.26 l=0.15
X14 a_74152_n2624# a_73934_n2624# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X15 a_80522_n2634# a_74152_n2624# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X16 charge_pump1_2/clk_in a_106522_n2434# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X17 a_74152_n2624# a_73934_n2624# charge_pump1_2/vdd charge_pump1_2/vdd sky130_fd_pr__pfet_01v8 ad=0.365 pd=3.1 as=0.365 ps=3.1 w=1.26 l=0.15
X18 a_80522_n2634# a_74152_n2624# charge_pump1_2/vdd charge_pump1_2/vdd sky130_fd_pr__pfet_01v8 ad=0.365 pd=3.1 as=0.365 ps=3.1 w=1.26 l=0.15
X19 a_99934_n2424# charge_pump1_reverse_1/clock_1/clk_in VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X20 charge_pump1_2/clk_in a_106522_n2434# charge_pump1_2/vdd charge_pump1_2/vdd sky130_fd_pr__pfet_01v8 ad=0.365 pd=3.1 as=0.365 ps=3.1 w=1.26 l=0.15
X21 a_99934_n2424# charge_pump1_reverse_1/clock_1/clk_in charge_pump1_2/vdd charge_pump1_2/vdd sky130_fd_pr__pfet_01v8 ad=0.365 pd=3.1 as=0.365 ps=3.1 w=1.26 l=0.15
X22 a_100152_n2424# a_99934_n2424# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X23 a_73934_n2624# charge_pump1_1/clk_in VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
C0 charge_pump1_2/in5 VSUBS 3.86f
C1 charge_pump1_2/vdd charge_pump1_2/in5 3.75f
C2 charge_pump1_1/a_3340_18086# VSUBS 6.14f
C3 charge_pump1_2/in3 VSUBS 3.87f
C4 charge_pump1_2/vdd charge_pump1_reverse_0/clock_1/clk_in 4.85f
C5 charge_pump1_2/vdd charge_pump1_2/in3 3.75f
C6 charge_pump1_2/vdd VSUBS 30f
C7 VSUBS charge_pump1_2/in8 3.71f
C8 charge_pump1_2/in2 VSUBS 3.88f
C9 charge_pump1_2/vdd charge_pump1_2/in8 3.69f
C10 charge_pump1_2/in2 charge_pump1_2/vdd 3.75f
C11 charge_pump1_1/clk_in charge_pump1_2/vdd 5.6f
C12 charge_pump1_2/in7 VSUBS 3.79f
C13 charge_pump1_2/clk_in charge_pump1_2/vdd 2.83f
C14 charge_pump1_2/vdd charge_pump1_2/in7 3.66f
C15 charge_pump1_2/in1 VSUBS 3.7f
C16 charge_pump1_2/in6 VSUBS 3.91f
C17 VSUBS charge_pump1_2/a_3340_18086# 6.04f
C18 charge_pump1_2/in1 charge_pump1_2/vdd 3.69f
C19 charge_pump1_2/vdd charge_pump1_reverse_1/clock_1/clk_in 5.61f
C20 charge_pump1_0/clk_in charge_pump1_2/vdd 4.6f
C21 charge_pump1_2/vdd charge_pump1_2/in6 3.78f
C22 charge_pump1_2/in4 VSUBS 3.86f
C23 charge_pump1_2/vdd charge_pump1_2/in4 3.75f
C24 charge_pump1_reverse_1/input1 0 22.9f
C25 charge_pump1_reverse_1/input2 0 22.4f
C26 charge_pump1_reverse_1/capacitors_1_12/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C27 charge_pump1_reverse_1/capacitors_1_12/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C28 charge_pump1_reverse_1/capacitors_1_12/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 0 2.66f
C29 charge_pump1_reverse_1/capacitors_1_13/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C30 charge_pump1_reverse_1/capacitors_1_13/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C31 charge_pump1_reverse_1/capacitors_1_13/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 0 2.66f
C32 charge_pump1_reverse_1/capacitors_1_11/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C33 charge_pump1_reverse_1/capacitors_1_11/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C34 charge_pump1_reverse_1/capacitors_1_11/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 0 2.66f
C35 charge_pump1_reverse_1/capacitors_1_10/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C36 charge_pump1_reverse_1/capacitors_1_10/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C37 charge_pump1_reverse_1/capacitors_1_10/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 0 2.66f
C38 charge_pump1_reverse_1/m1_4341_n519# 0 3.86f
C39 charge_pump1_reverse_1/m1_12659_300# 0 2.73f
C40 charge_pump1_2/nmos_dnw3_0/vs 0 15.1f
C41 charge_pump1_reverse_1/capacitors_1_9/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C42 charge_pump1_reverse_1/capacitors_1_9/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C43 charge_pump1_reverse_1/capacitors_1_9/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 0 2.66f
C44 charge_pump1_reverse_1/capacitors_1_8/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C45 charge_pump1_reverse_1/capacitors_1_8/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C46 charge_pump1_reverse_1/capacitors_1_8/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 0 2.66f
C47 charge_pump1_reverse_1/capacitors_1_7/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C48 charge_pump1_reverse_1/capacitors_1_7/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C49 charge_pump1_reverse_1/capacitors_1_7/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 0 2.66f
C50 charge_pump1_reverse_1/capacitors_1_6/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C51 charge_pump1_reverse_1/capacitors_1_6/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C52 charge_pump1_reverse_1/capacitors_1_6/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 0 2.66f
C53 charge_pump1_reverse_1/capacitors_1_5/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C54 charge_pump1_reverse_1/capacitors_1_5/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C55 charge_pump1_reverse_1/capacitors_1_5/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 0 2.66f
C56 charge_pump1_reverse_1/capacitors_1_4/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C57 charge_pump1_reverse_1/capacitors_1_4/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C58 charge_pump1_reverse_1/capacitors_1_4/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 0 2.66f
C59 charge_pump1_reverse_1/capacitors_1_3/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C60 charge_pump1_reverse_1/capacitors_1_3/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C61 charge_pump1_reverse_1/capacitors_1_3/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 0 2.66f
C62 charge_pump1_reverse_1/capacitors_1_2/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C63 charge_pump1_reverse_1/capacitors_1_2/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C64 charge_pump1_reverse_1/capacitors_1_2/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 0 2.66f
C65 charge_pump1_reverse_1/capacitors_1_1/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C66 charge_pump1_reverse_1/capacitors_1_1/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C67 charge_pump1_reverse_1/capacitors_1_1/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 0 2.66f
C68 charge_pump1_reverse_1/capacitors_1_0/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C69 charge_pump1_reverse_1/capacitors_1_0/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C70 charge_pump1_reverse_1/capacitors_1_0/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 0 2.66f
C71 charge_pump1_2/in8 0 7.62f
C72 charge_pump1_reverse_1/capacitor_8_1/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C73 charge_pump1_reverse_1/clock_1/clk 0 88.1f
C74 charge_pump1_reverse_1/capacitor_8_1/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C75 charge_pump1_reverse_1/capacitor_8_1/capacitor_7_0/buffer_and_gate_0/in1 0 2.66f
C76 charge_pump1_reverse_1/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C77 charge_pump1_reverse_1/clock_1/clkb 0 96.8f
C78 charge_pump1_reverse_1/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C79 charge_pump1_reverse_1/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 0 2.66f
C80 charge_pump1_reverse_1/clock_1/a_2432_n962# 0 8.68f **FLOATING
C81 charge_pump1_reverse_1/clock_1/a_2020_n482# 0 2.57f **FLOATING
C82 charge_pump1_reverse_1/clock_1/a_344_102# 0 2.81f
C83 charge_pump1_reverse_1/clock_1/a_2402_572# 0 2.17f
C84 charge_pump1_reverse_1/clock_1/a_344_n986# 0 2.38f
C85 charge_pump1_reverse_1/clock_1/clk_in 0 14.7f
C86 charge_pump1_reverse_1/clock_1/a_3246_118# 0 6.83f
C87 charge_pump1_reverse_1/nmos_dnw3_0/clkb 0 2.01f
C88 charge_pump1_reverse_0/input1 0 22.9f
C89 charge_pump1_reverse_0/input2 0 22.4f
C90 charge_pump1_reverse_0/capacitors_1_12/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C91 charge_pump1_reverse_0/capacitors_1_12/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C92 charge_pump1_reverse_0/capacitors_1_12/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 0 2.66f
C93 charge_pump1_reverse_0/capacitors_1_13/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C94 charge_pump1_reverse_0/capacitors_1_13/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C95 charge_pump1_reverse_0/capacitors_1_13/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 0 2.66f
C96 charge_pump1_reverse_0/capacitors_1_11/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C97 charge_pump1_reverse_0/capacitors_1_11/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C98 charge_pump1_reverse_0/capacitors_1_11/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 0 2.66f
C99 charge_pump1_reverse_0/capacitors_1_10/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C100 charge_pump1_reverse_0/capacitors_1_10/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C101 charge_pump1_reverse_0/capacitors_1_10/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 0 2.66f
C102 charge_pump1_reverse_0/m1_4341_n519# 0 3.86f
C103 charge_pump1_reverse_0/m1_12659_300# 0 2.73f
C104 charge_pump1_1/nmos_dnw3_0/vs 0 15.1f
C105 charge_pump1_reverse_0/capacitors_1_9/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C106 charge_pump1_reverse_0/capacitors_1_9/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C107 charge_pump1_reverse_0/capacitors_1_9/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 0 2.66f
C108 charge_pump1_reverse_0/capacitors_1_8/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C109 charge_pump1_reverse_0/capacitors_1_8/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C110 charge_pump1_reverse_0/capacitors_1_8/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 0 2.66f
C111 charge_pump1_reverse_0/capacitors_1_7/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C112 charge_pump1_reverse_0/capacitors_1_7/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C113 charge_pump1_reverse_0/capacitors_1_7/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 0 2.66f
C114 charge_pump1_reverse_0/capacitors_1_6/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C115 charge_pump1_reverse_0/capacitors_1_6/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C116 charge_pump1_reverse_0/capacitors_1_6/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 0 2.66f
C117 charge_pump1_reverse_0/capacitors_1_5/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C118 charge_pump1_reverse_0/capacitors_1_5/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C119 charge_pump1_reverse_0/capacitors_1_5/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 0 2.66f
C120 charge_pump1_reverse_0/capacitors_1_4/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C121 charge_pump1_reverse_0/capacitors_1_4/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C122 charge_pump1_reverse_0/capacitors_1_4/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 0 2.66f
C123 charge_pump1_reverse_0/capacitors_1_3/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C124 charge_pump1_reverse_0/capacitors_1_3/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C125 charge_pump1_reverse_0/capacitors_1_3/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 0 2.66f
C126 charge_pump1_reverse_0/capacitors_1_2/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C127 charge_pump1_reverse_0/capacitors_1_2/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C128 charge_pump1_reverse_0/capacitors_1_2/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 0 2.66f
C129 charge_pump1_reverse_0/capacitors_1_1/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C130 charge_pump1_reverse_0/capacitors_1_1/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C131 charge_pump1_reverse_0/capacitors_1_1/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 0 2.66f
C132 charge_pump1_reverse_0/capacitors_1_0/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C133 charge_pump1_reverse_0/capacitors_1_0/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C134 charge_pump1_reverse_0/capacitors_1_0/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 0 2.66f
C135 charge_pump1_reverse_0/capacitor_8_1/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C136 charge_pump1_reverse_0/clock_1/clk 0 88.1f
C137 charge_pump1_reverse_0/capacitor_8_1/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C138 charge_pump1_reverse_0/capacitor_8_1/capacitor_7_0/buffer_and_gate_0/in1 0 2.66f
C139 VSUBS 0 0.35p
C140 charge_pump1_reverse_0/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C141 charge_pump1_reverse_0/clock_1/clkb 0 96.8f
C142 charge_pump1_reverse_0/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C143 charge_pump1_reverse_0/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 0 2.66f
C144 charge_pump1_reverse_0/clock_1/a_2432_n962# 0 8.68f **FLOATING
C145 charge_pump1_reverse_0/clock_1/a_2020_n482# 0 2.57f **FLOATING
C146 charge_pump1_reverse_0/clock_1/a_344_102# 0 2.81f
C147 charge_pump1_reverse_0/clock_1/a_2402_572# 0 2.17f
C148 charge_pump1_reverse_0/clock_1/a_344_n986# 0 2.38f
C149 charge_pump1_reverse_0/clock_1/clk_in 0 12.2f
C150 charge_pump1_reverse_0/clock_1/a_3246_118# 0 6.83f
C151 charge_pump1_reverse_0/nmos_dnw3_0/clkb 0 2.01f
C152 charge_pump1_2/input1 0 22.5f
C153 charge_pump1_2/input2 0 22.2f
C154 charge_pump1_2/capacitors_1_12/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C155 charge_pump1_2/capacitors_1_12/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C156 charge_pump1_2/capacitors_1_12/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 0 2.66f
C157 charge_pump1_2/capacitors_1_13/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C158 charge_pump1_2/capacitors_1_13/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C159 charge_pump1_2/capacitors_1_13/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 0 2.66f
C160 charge_pump1_2/capacitors_1_11/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C161 charge_pump1_2/capacitors_1_11/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C162 charge_pump1_2/capacitors_1_11/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 0 2.66f
C163 charge_pump1_2/capacitors_1_10/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C164 charge_pump1_2/capacitors_1_10/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C165 charge_pump1_2/capacitors_1_10/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 0 2.66f
C166 charge_pump1_2/m1_4341_n519# 0 3.77f
C167 charge_pump1_2/m1_12659_300# 0 2.54f
C168 charge_pump1_2/m1_12464_n576# 0 4.25f
C169 charge_pump1_2/capacitors_1_9/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C170 charge_pump1_2/capacitors_1_9/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C171 charge_pump1_2/capacitors_1_9/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 0 2.66f
C172 charge_pump1_2/capacitors_1_8/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C173 charge_pump1_2/capacitors_1_8/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C174 charge_pump1_2/capacitors_1_8/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 0 2.66f
C175 charge_pump1_2/capacitors_1_7/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C176 charge_pump1_2/capacitors_1_7/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C177 charge_pump1_2/capacitors_1_7/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 0 2.66f
C178 charge_pump1_2/capacitors_1_6/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C179 charge_pump1_2/capacitors_1_6/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C180 charge_pump1_2/capacitors_1_6/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 0 2.66f
C181 charge_pump1_2/capacitors_1_5/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C182 charge_pump1_2/capacitors_1_5/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C183 charge_pump1_2/capacitors_1_5/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 0 2.66f
C184 charge_pump1_2/capacitors_1_4/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C185 charge_pump1_2/capacitors_1_4/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C186 charge_pump1_2/capacitors_1_4/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 0 2.66f
C187 charge_pump1_2/capacitors_1_3/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C188 charge_pump1_2/capacitors_1_3/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C189 charge_pump1_2/capacitors_1_3/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 0 2.66f
C190 charge_pump1_2/capacitors_1_2/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C191 charge_pump1_2/capacitors_1_2/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C192 charge_pump1_2/capacitors_1_2/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 0 2.66f
C193 charge_pump1_2/capacitors_1_1/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C194 charge_pump1_2/capacitors_1_1/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C195 charge_pump1_2/capacitors_1_1/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 0 2.66f
C196 charge_pump1_2/capacitors_1_0/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C197 charge_pump1_2/capacitors_1_0/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C198 charge_pump1_2/capacitors_1_0/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 0 2.66f
C199 charge_pump1_2/capacitor_8_1/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C200 charge_pump1_2/clock_0/clkb 0 86.1f
C201 charge_pump1_2/capacitor_8_1/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C202 charge_pump1_2/capacitor_8_1/capacitor_7_0/buffer_and_gate_0/in1 0 2.66f
C203 charge_pump1_2/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C204 charge_pump1_2/clock_0/clk 0 85.5f
C205 charge_pump1_2/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C206 charge_pump1_2/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 0 2.66f
C207 charge_pump1_2/clock_0/a_2432_n962# 0 8.68f **FLOATING
C208 charge_pump1_2/clock_0/a_2020_n482# 0 2.57f **FLOATING
C209 charge_pump1_2/clock_0/a_344_102# 0 2.81f
C210 charge_pump1_2/clock_0/a_2402_572# 0 2.17f
C211 charge_pump1_2/clock_0/a_344_n986# 0 2.38f
C212 charge_pump1_2/clk_in 0 11.3f
C213 charge_pump1_2/clock_0/a_3246_118# 0 6.83f
C214 charge_pump1_2/nmos_dnw3_0/clkb 0 2.34f
C215 charge_pump1_1/input1 0 22.5f
C216 charge_pump1_1/input2 0 22.2f
C217 charge_pump1_1/capacitors_1_12/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C218 charge_pump1_1/capacitors_1_12/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C219 charge_pump1_1/capacitors_1_12/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 0 2.66f
C220 charge_pump1_1/capacitors_1_13/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C221 charge_pump1_1/capacitors_1_13/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C222 charge_pump1_1/capacitors_1_13/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 0 2.66f
C223 charge_pump1_1/capacitors_1_11/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C224 charge_pump1_1/capacitors_1_11/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C225 charge_pump1_1/capacitors_1_11/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 0 2.66f
C226 charge_pump1_1/capacitors_1_10/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C227 charge_pump1_1/capacitors_1_10/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C228 charge_pump1_1/capacitors_1_10/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 0 2.66f
C229 charge_pump1_1/m1_4341_n519# 0 3.77f
C230 charge_pump1_1/m1_12659_300# 0 2.54f
C231 charge_pump1_reverse_1/nmos_dnw3_0/vs 0 14.5f
C232 charge_pump1_1/capacitors_1_9/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C233 charge_pump1_1/capacitors_1_9/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C234 charge_pump1_1/capacitors_1_9/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 0 2.66f
C235 charge_pump1_2/in7 0 7.2f
C236 charge_pump1_1/capacitors_1_8/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C237 charge_pump1_1/capacitors_1_8/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C238 charge_pump1_1/capacitors_1_8/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 0 2.66f
C239 charge_pump1_2/in6 0 7.22f
C240 charge_pump1_1/capacitors_1_7/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C241 charge_pump1_1/capacitors_1_7/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C242 charge_pump1_1/capacitors_1_7/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 0 2.66f
C243 charge_pump1_2/in5 0 7.33f
C244 charge_pump1_1/capacitors_1_6/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C245 charge_pump1_1/capacitors_1_6/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C246 charge_pump1_1/capacitors_1_6/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 0 2.66f
C247 charge_pump1_1/capacitors_1_5/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C248 charge_pump1_1/capacitors_1_5/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C249 charge_pump1_1/capacitors_1_5/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 0 2.66f
C250 charge_pump1_1/capacitors_1_4/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C251 charge_pump1_1/capacitors_1_4/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C252 charge_pump1_1/capacitors_1_4/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 0 2.66f
C253 charge_pump1_1/capacitors_1_3/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C254 charge_pump1_1/capacitors_1_3/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C255 charge_pump1_1/capacitors_1_3/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 0 2.66f
C256 charge_pump1_2/in3 0 7.21f
C257 charge_pump1_1/capacitors_1_2/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C258 charge_pump1_1/capacitors_1_2/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C259 charge_pump1_1/capacitors_1_2/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 0 2.66f
C260 charge_pump1_2/in2 0 7.21f
C261 charge_pump1_1/capacitors_1_1/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C262 charge_pump1_1/capacitors_1_1/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C263 charge_pump1_1/capacitors_1_1/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 0 2.66f
C264 charge_pump1_1/capacitors_1_0/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C265 charge_pump1_1/capacitors_1_0/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C266 charge_pump1_1/capacitors_1_0/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 0 2.66f
C267 charge_pump1_2/in1 0 6.91f
C268 charge_pump1_1/capacitor_8_1/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C269 charge_pump1_1/clock_0/clkb 0 86.1f
C270 charge_pump1_1/capacitor_8_1/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C271 charge_pump1_1/capacitor_8_1/capacitor_7_0/buffer_and_gate_0/in1 0 2.66f
C272 charge_pump1_1/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C273 charge_pump1_1/clock_0/clk 0 85.5f
C274 charge_pump1_1/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C275 charge_pump1_1/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 0 2.66f
C276 charge_pump1_1/clock_0/a_2432_n962# 0 8.68f **FLOATING
C277 charge_pump1_1/clock_0/a_2020_n482# 0 2.57f **FLOATING
C278 charge_pump1_1/clock_0/a_344_102# 0 2.81f
C279 charge_pump1_1/clock_0/a_2402_572# 0 2.17f
C280 charge_pump1_1/clock_0/a_344_n986# 0 2.38f
C281 charge_pump1_1/clk_in 0 18.2f
C282 charge_pump1_1/clock_0/a_3246_118# 0 6.83f
C283 charge_pump1_1/nmos_dnw3_0/clkb 0 2.34f
C284 charge_pump1_0/input1 0 22.5f
C285 charge_pump1_0/input2 0 22.2f
C286 charge_pump1_0/capacitors_1_12/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C287 charge_pump1_0/capacitors_1_12/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C288 charge_pump1_0/capacitors_1_12/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 0 2.66f
C289 charge_pump1_0/capacitors_1_13/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C290 charge_pump1_0/capacitors_1_13/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C291 charge_pump1_0/capacitors_1_13/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 0 2.66f
C292 charge_pump1_0/capacitors_1_11/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C293 charge_pump1_0/capacitors_1_11/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C294 charge_pump1_0/capacitors_1_11/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 0 2.66f
C295 charge_pump1_0/capacitors_1_10/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C296 charge_pump1_0/capacitors_1_10/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C297 charge_pump1_0/capacitors_1_10/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 0 2.66f
C298 charge_pump1_0/m1_4341_n519# 0 3.77f
C299 charge_pump1_0/m1_12659_300# 0 2.54f
C300 charge_pump1_reverse_0/nmos_dnw3_0/vs 0 14.7f
C301 charge_pump1_0/capacitors_1_9/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C302 charge_pump1_0/capacitors_1_9/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C303 charge_pump1_0/capacitors_1_9/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 0 2.66f
C304 charge_pump1_0/capacitors_1_8/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C305 charge_pump1_0/capacitors_1_8/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C306 charge_pump1_0/capacitors_1_8/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 0 2.66f
C307 charge_pump1_0/capacitors_1_7/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C308 charge_pump1_0/capacitors_1_7/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C309 charge_pump1_0/capacitors_1_7/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 0 2.66f
C310 charge_pump1_0/capacitors_1_6/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C311 charge_pump1_0/capacitors_1_6/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C312 charge_pump1_0/capacitors_1_6/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 0 2.66f
C313 charge_pump1_2/in4 0 7.33f
C314 charge_pump1_0/capacitors_1_5/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C315 charge_pump1_0/capacitors_1_5/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C316 charge_pump1_0/capacitors_1_5/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 0 2.66f
C317 charge_pump1_0/capacitors_1_4/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C318 charge_pump1_0/capacitors_1_4/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C319 charge_pump1_0/capacitors_1_4/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 0 2.66f
C320 charge_pump1_0/capacitors_1_3/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C321 charge_pump1_0/capacitors_1_3/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C322 charge_pump1_0/capacitors_1_3/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 0 2.66f
C323 charge_pump1_0/capacitors_1_2/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C324 charge_pump1_0/capacitors_1_2/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C325 charge_pump1_0/capacitors_1_2/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 0 2.66f
C326 charge_pump1_0/capacitors_1_1/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C327 charge_pump1_0/capacitors_1_1/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C328 charge_pump1_0/capacitors_1_1/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 0 2.66f
C329 charge_pump1_0/capacitors_1_0/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C330 charge_pump1_0/capacitors_1_0/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C331 charge_pump1_0/capacitors_1_0/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 0 2.66f
C332 charge_pump1_0/capacitor_8_1/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C333 charge_pump1_0/clock_0/clkb 0 86.1f
C334 charge_pump1_0/capacitor_8_1/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C335 charge_pump1_0/capacitor_8_1/capacitor_7_0/buffer_and_gate_0/in1 0 2.66f
C336 charge_pump1_0/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C337 charge_pump1_0/clock_0/clk 0 85.5f
C338 charge_pump1_0/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C339 charge_pump1_2/vdd 0 2.37p
C340 charge_pump1_0/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 0 2.66f
C341 charge_pump1_0/clock_0/a_2432_n962# 0 8.68f **FLOATING
C342 charge_pump1_0/clock_0/a_2020_n482# 0 2.57f **FLOATING
C343 charge_pump1_0/clock_0/a_344_102# 0 2.81f
C344 charge_pump1_0/clock_0/a_2402_572# 0 2.17f
C345 charge_pump1_0/clock_0/a_344_n986# 0 2.38f
C346 charge_pump1_0/clk_in 0 21f
C347 charge_pump1_0/clock_0/a_3246_118# 0 6.83f
C348 charge_pump1_0/nmos_dnw3_0/clkb 0 2.34f
C349 charge_pump1_0/nmos_dnw3_0/vs 0 10.4f
.ends

.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
X0 VPWR VGND VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0.452 ps=4.52 w=0.87 l=0.59
X1 VGND VPWR VGND VNB sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0.286 ps=3.24 w=0.55 l=0.59
.ends

.subckt sky130_fd_sc_hd__a21oi_1 A1 A2 B1 VGND VNB VPB VPWR Y
X0 a_199_47# A1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.0959 pd=0.945 as=0.091 ps=0.93 w=0.65 l=0.15
X1 a_113_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.147 ps=1.29 w=1 l=0.15
X2 Y B1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.172 ps=1.83 w=0.65 l=0.15
X3 VPWR A1 a_113_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.147 pd=1.29 as=0.14 ps=1.28 w=1 l=0.15
X4 a_113_297# B1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X5 VGND A2 a_199_47# VNB sky130_fd_pr__nfet_01v8 ad=0.172 pd=1.83 as=0.0959 ps=0.945 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__o31a_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
X0 a_103_199# B1 a_253_47# VNB sky130_fd_pr__nfet_01v8 ad=0.201 pd=1.92 as=0.107 ps=0.98 w=0.65 l=0.15
X1 VPWR a_103_199# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=1.39 as=0.36 ps=2.72 w=1 l=0.15
X2 a_337_297# A2 a_253_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.135 ps=1.27 w=1 l=0.15
X3 a_103_199# A3 a_337_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.213 pd=1.42 as=0.165 ps=1.33 w=1 l=0.15
X4 a_253_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.195 ps=1.39 w=1 l=0.15
X5 VPWR B1 a_103_199# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.345 pd=2.69 as=0.213 ps=1.42 w=1 l=0.15
X6 VGND a_103_199# X VNB sky130_fd_pr__nfet_01v8 ad=0.127 pd=1.04 as=0.234 ps=2.02 w=0.65 l=0.15
X7 a_253_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.127 ps=1.04 w=0.65 l=0.15
X8 a_253_47# A3 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.107 ps=0.98 w=0.65 l=0.15
X9 VGND A2 a_253_47# VNB sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.0878 ps=0.92 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
X0 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X1 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.149 ps=1.33 w=1 l=0.15
X2 VPWR A a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.33 as=0.166 ps=1.8 w=0.64 l=0.15
X3 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X4 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.172 pd=1.83 as=0.0878 ps=0.92 w=0.65 l=0.15
X5 VGND A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__or3_1 A B C VGND VNB VPB VPWR X
X0 X a_29_53# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.148 ps=1.34 w=1 l=0.15
X1 a_111_297# C a_29_53# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.109 ps=1.36 w=0.42 l=0.15
X2 X a_29_53# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.102 ps=0.99 w=0.65 l=0.15
X3 a_183_297# B a_111_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X4 VPWR A a_183_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.148 pd=1.34 as=0.0693 ps=0.75 w=0.42 l=0.15
X5 a_29_53# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X6 VGND C a_29_53# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X7 VGND A a_29_53# VNB sky130_fd_pr__nfet_01v8 ad=0.102 pd=0.99 as=0.0567 ps=0.69 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__clkbuf_4 A VGND VNB VPB VPWR X
X0 VPWR A a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.265 ps=2.53 w=1 l=0.15
X1 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0588 ps=0.7 w=0.42 l=0.15
X2 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X5 VGND A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0703 pd=0.755 as=0.111 ps=1.37 w=0.42 l=0.15
X6 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.14 ps=1.28 w=1 l=0.15
X7 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0703 ps=0.755 w=0.42 l=0.15
X8 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.165 ps=1.33 w=1 l=0.15
X9 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
.ends

.subckt sky130_fd_sc_hd__o21a_1 A1 A2 B1 VGND VNB VPB VPWR X
X0 VPWR A1 a_382_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.153 ps=1.3 w=1 l=0.15
X1 a_297_47# B1 a_79_21# VNB sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.96 as=0.169 ps=1.82 w=0.65 l=0.15
X2 a_297_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X3 VGND A2 a_297_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.101 ps=0.96 w=0.65 l=0.15
X4 VPWR a_79_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.327 pd=1.65 as=0.28 ps=2.56 w=1 l=0.15
X5 a_79_21# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=1.39 as=0.327 ps=1.65 w=1 l=0.15
X6 a_382_297# A2 a_79_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.153 pd=1.3 as=0.195 ps=1.39 w=1 l=0.15
X7 VGND a_79_21# X VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
X0 VPWR VGND VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0.452 ps=4.52 w=0.87 l=2.89
X1 VGND VPWR VGND VNB sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0.286 ps=3.24 w=0.55 l=2.89
.ends

.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
X0 VPWR VGND VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0.452 ps=4.52 w=0.87 l=1.97
X1 VGND VPWR VGND VNB sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0.286 ps=3.24 w=0.55 l=1.97
.ends

.subckt sky130_fd_sc_hd__nor3b_1 A B C_N VGND VNB VPB VPWR Y
X0 VGND a_91_199# Y VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.221 ps=1.98 w=0.65 l=0.15
X1 Y B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X2 VPWR A a_245_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.146 pd=1.34 as=0.135 ps=1.27 w=1 l=0.15
X3 a_91_199# C_N VGND VNB sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.1 ps=0.985 w=0.42 l=0.15
X4 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.985 as=0.0878 ps=0.92 w=0.65 l=0.15
X5 a_245_297# B a_161_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6 a_91_199# C_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.146 ps=1.34 w=0.42 l=0.15
X7 a_161_297# a_91_199# Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.32 ps=2.64 w=1 l=0.15
.ends

.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
X0 VPWR VGND VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0.452 ps=4.52 w=0.87 l=1.05
X1 VGND VPWR VGND VNB sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0.286 ps=3.24 w=0.55 l=1.05
.ends

.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
X0 VPWR A a_110_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X5 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X6 a_110_47# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X7 a_110_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X8 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X9 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X10 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X11 a_110_47# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X12 VGND A a_110_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X13 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.0578 pd=0.695 as=0.0588 ps=0.7 w=0.42 l=0.15
X14 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X15 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X16 VGND A a_110_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X17 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.111 pd=1.37 as=0.0588 ps=0.7 w=0.42 l=0.15
X18 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.138 pd=1.27 as=0.14 ps=1.28 w=1 l=0.15
X19 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X20 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.138 ps=1.27 w=1 l=0.15
X21 a_110_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.111 ps=1.37 w=0.42 l=0.15
X22 VPWR A a_110_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X23 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X24 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X25 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X26 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X27 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X28 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X29 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X30 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X31 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X32 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X33 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X34 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X35 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X36 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X37 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X38 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X39 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0578 ps=0.695 w=0.42 l=0.15
.ends

.subckt sky130_ef_sc_hd__decap_12 VGND VPWR VPB VNB
X0 VPWR VGND VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0.452 ps=4.52 w=0.87 l=4.73
X1 VGND VPWR VGND VNB sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0.286 ps=3.24 w=0.55 l=4.73
.ends

.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
X0 VPWR A a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.162 pd=1.33 as=0.265 ps=2.53 w=1 l=0.15
X1 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2 VGND A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0683 pd=0.745 as=0.111 ps=1.37 w=0.42 l=0.15
X3 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.162 ps=1.33 w=1 l=0.15
X4 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0683 ps=0.745 w=0.42 l=0.15
X5 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
X0 VPWR a_75_212# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X1 a_75_212# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X2 a_75_212# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X3 VGND a_75_212# X VNB sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
.ends

.subckt sky130_fd_sc_hd__dlymetal6s2s_1 A VGND VNB VPB VPWR X
X0 a_558_47# a_381_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.141 ps=1.33 w=1 l=0.15
X1 VGND X a_381_47# VNB sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X2 a_841_47# a_664_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.141 ps=1.33 w=1 l=0.15
X3 VPWR A a_62_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.141 pd=1.33 as=0.109 ps=1.36 w=0.42 l=0.15
X4 VGND A a_62_47# VNB sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X5 a_558_47# a_381_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X6 X a_62_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.141 ps=1.33 w=1 l=0.15
X7 VPWR X a_381_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.141 pd=1.33 as=0.109 ps=1.36 w=0.42 l=0.15
X8 a_841_47# a_664_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X9 X a_62_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X10 VPWR a_558_47# a_664_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.141 pd=1.33 as=0.109 ps=1.36 w=0.42 l=0.15
X11 VGND a_558_47# a_664_47# VNB sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__dfrtp_1 CLK D RESET_B VGND VNB VPB VPWR Q
X0 a_1217_47# a_27_47# a_1108_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X1 a_805_47# a_761_289# a_639_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.14 ps=1.1 w=0.42 l=0.15
X2 a_1108_47# a_193_47# a_761_289# VNB sky130_fd_pr__nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X3 a_1283_21# a_1108_47# a_1462_47# VNB sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.064 ps=0.725 w=0.42 l=0.15
X4 a_651_413# a_27_47# a_543_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.116 pd=0.97 as=0.0724 ps=0.765 w=0.42 l=0.15
X5 VGND RESET_B a_805_47# VNB sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X6 Q a_1283_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.301 ps=2.66 w=1 l=0.15
X7 VPWR CLK a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X8 a_448_47# D VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.109 ps=1.36 w=0.42 l=0.15
X9 a_761_289# a_543_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.135 ps=1.15 w=0.64 l=0.15
X10 a_193_47# a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X11 a_1108_47# a_27_47# a_761_289# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.129 ps=1.18 w=0.42 l=0.15
X12 a_543_47# a_27_47# a_448_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X13 a_1462_47# RESET_B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.064 pd=0.725 as=0.125 ps=1.01 w=0.42 l=0.15
X14 a_543_47# a_193_47# a_448_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0724 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X15 a_448_47# D VGND VNB sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.221 ps=1.89 w=0.42 l=0.15
X16 VPWR a_1283_21# a_1270_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X17 VPWR a_1108_47# a_1283_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.113 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X18 a_1270_413# a_193_47# a_1108_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X19 a_193_47# a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X20 a_1283_21# RESET_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X21 VPWR a_761_289# a_651_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0703 pd=0.755 as=0.116 ps=0.97 w=0.42 l=0.15
X22 Q a_1283_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.209 ps=2.02 w=0.65 l=0.15
X23 a_639_47# a_193_47# a_543_47# VNB sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X24 VGND a_1283_21# a_1217_47# VNB sky130_fd_pr__nfet_01v8 ad=0.125 pd=1.01 as=0.0669 ps=0.75 w=0.42 l=0.15
X25 a_651_413# RESET_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0703 ps=0.755 w=0.42 l=0.15
X26 VGND CLK a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X27 a_761_289# a_543_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.129 pd=1.18 as=0.218 ps=2.2 w=0.84 l=0.15
.ends

.subckt sky130_fd_sc_hd__and2_1 A B VGND VNB VPB VPWR X
X0 VPWR B a_59_75# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.167 pd=1.39 as=0.0567 ps=0.69 w=0.42 l=0.15
X1 X a_59_75# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.475 pd=2.95 as=0.167 ps=1.39 w=1 l=0.15
X2 VGND B a_145_75# VNB sky130_fd_pr__nfet_01v8 ad=0.112 pd=1.04 as=0.0567 ps=0.69 w=0.42 l=0.15
X3 a_59_75# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.118 ps=1.4 w=0.42 l=0.15
X4 X a_59_75# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.112 ps=1.04 w=0.65 l=0.15
X5 a_145_75# A a_59_75# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.118 ps=1.4 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__dlygate4sd3_1 A VGND VNB VPB VPWR X
X0 VPWR A a_49_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X1 VGND a_285_47# a_391_47# VNB sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.5
X2 X a_391_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.141 ps=1.33 w=1 l=0.15
X3 VGND A a_49_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X4 VPWR a_285_47# a_391_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.141 pd=1.33 as=0.109 ps=1.36 w=0.42 l=0.5
X5 a_285_47# a_49_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.5
X6 a_285_47# a_49_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.5
X7 X a_391_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__nor2_2 A B VGND VNB VPB VPWR Y
X0 Y B a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1 Y B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X2 a_27_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X4 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.182 ps=1.86 w=0.65 l=0.15
X5 VGND B Y VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X6 VPWR A a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=2.56 w=1 l=0.15
X7 a_27_297# B Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
.ends

.subckt sky130_fd_sc_hd__o32a_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
X0 a_77_199# B2 a_227_47# VNB sky130_fd_pr__nfet_01v8 ad=0.133 pd=1.06 as=0.127 ps=1.04 w=0.65 l=0.15
X1 a_323_297# A2 a_227_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=1.39 as=0.165 ps=1.33 w=1 l=0.15
X2 a_227_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.135 ps=1.27 w=1 l=0.15
X3 a_227_47# B1 a_77_199# VNB sky130_fd_pr__nfet_01v8 ad=0.189 pd=1.88 as=0.133 ps=1.06 w=0.65 l=0.15
X4 VGND a_77_199# X VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5 VPWR B1 a_539_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.205 ps=1.41 w=1 l=0.15
X6 a_227_47# A3 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.127 pd=1.04 as=0.127 ps=1.04 w=0.65 l=0.15
X7 VPWR a_77_199# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.335 ps=2.67 w=1 l=0.15
X8 a_77_199# A3 a_323_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=1.39 as=0.195 ps=1.39 w=1 l=0.15
X9 VGND A2 a_227_47# VNB sky130_fd_pr__nfet_01v8 ad=0.127 pd=1.04 as=0.107 ps=0.98 w=0.65 l=0.15
X10 a_227_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.0878 ps=0.92 w=0.65 l=0.15
X11 a_539_297# B2 a_77_199# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=1.41 as=0.195 ps=1.39 w=1 l=0.15
.ends

.subckt scanchain VDD data_out[0] data_out[1] data_out[2] data_out[3] data_out[4]
+ data_out[5] data_out[6] data_out[7] scan_out GND
XPHY_EDGE_ROW_0_Left_12 GND GND VDD VDD sky130_fd_sc_hd__decap_3
X_66_ net1 _09_ _08_ GND GND VDD VDD _33_ sky130_fd_sc_hd__a21oi_1
X_49_ _11_ _18_ _19_ _20_ GND GND VDD VDD _02_ sky130_fd_sc_hd__o31a_1
Xoutput7 net7 GND GND VDD VDD data_out[1] sky130_fd_sc_hd__buf_2
X_65_ _11_ _30_ _31_ _32_ GND GND VDD VDD _06_ sky130_fd_sc_hd__o31a_1
XFILLER_0_9_39 GND GND VDD VDD sky130_fd_sc_hd__decap_3
X_48_ _12_ net1 net17 GND GND VDD VDD _20_ sky130_fd_sc_hd__or3_1
XPHY_EDGE_ROW_6_Right_6 GND GND VDD VDD sky130_fd_sc_hd__decap_3
Xoutput10 net10 GND GND VDD VDD data_out[4] sky130_fd_sc_hd__clkbuf_4
Xoutput8 net8 GND GND VDD VDD data_out[2] sky130_fd_sc_hd__buf_2
X_64_ net3 net1 net18 GND GND VDD VDD _32_ sky130_fd_sc_hd__or3_1
X_47_ _12_ _09_ net7 GND GND VDD VDD _19_ sky130_fd_sc_hd__o21a_1
XFILLER_0_9_3 GND GND VDD VDD sky130_fd_sc_hd__decap_8
Xoutput11 net11 GND GND VDD VDD data_out[5] sky130_fd_sc_hd__buf_2
Xoutput9 net9 GND GND VDD VDD data_out[3] sky130_fd_sc_hd__buf_2
X_63_ _12_ net5 net11 GND GND VDD VDD _31_ sky130_fd_sc_hd__o21a_1
XFILLER_0_10_22 GND GND VDD VDD sky130_fd_sc_hd__decap_6
X_46_ _08_ _09_ net9 GND GND VDD VDD _18_ sky130_fd_sc_hd__nor3b_1
XPHY_EDGE_ROW_4_Left_16 GND GND VDD VDD sky130_fd_sc_hd__decap_3
Xoutput12 net12 GND GND VDD VDD data_out[6] sky130_fd_sc_hd__buf_2
X_62_ _08_ _09_ net13 GND GND VDD VDD _30_ sky130_fd_sc_hd__nor3b_1
X_45_ _11_ _15_ _16_ _17_ GND GND VDD VDD _01_ sky130_fd_sc_hd__o31a_1
Xoutput13 net13 GND GND VDD VDD data_out[7] sky130_fd_sc_hd__clkbuf_4
X_61_ _11_ _27_ _28_ _29_ GND GND VDD VDD _05_ sky130_fd_sc_hd__o31a_1
X_44_ _12_ net1 net7 GND GND VDD VDD _17_ sky130_fd_sc_hd__or3_1
Xoutput14 net14 GND GND VDD VDD scan_out sky130_fd_sc_hd__clkbuf_4
X_60_ net3 net1 net11 GND GND VDD VDD _29_ sky130_fd_sc_hd__or3_1
X_43_ _08_ _09_ net6 GND GND VDD VDD _16_ sky130_fd_sc_hd__o21a_1
XPHY_EDGE_ROW_1_Right_1 GND GND VDD VDD sky130_fd_sc_hd__decap_3
X_42_ _08_ _09_ net8 GND GND VDD VDD _15_ sky130_fd_sc_hd__nor3b_1
XPHY_EDGE_ROW_11_Left_23 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_0_1_13 GND GND VDD VDD sky130_fd_sc_hd__decap_4
Xclkbuf_0_clk clkbuf_0_clk/A GND GND VDD VDD clknet_0_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_4_24 GND GND VDD VDD sky130_fd_sc_hd__decap_4
X_41_ _10_ _11_ _13_ _14_ GND GND VDD VDD _00_ sky130_fd_sc_hd__o31a_1
XFILLER_0_7_46 GND GND VDD VDD sky130_fd_sc_hd__decap_8
X_40_ _12_ net1 net6 GND GND VDD VDD _14_ sky130_fd_sc_hd__or3_1
XPHY_EDGE_ROW_5_Right_5 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_0_7_7 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_10_29 GND GND VDD VDD sky130_fd_sc_hd__decap_8
XFILLER_0_1_38 GND GND VDD VDD sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_11_Right_11 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_0_7_37 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_3_Left_15 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_0_5_6 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_0_11_41 GND VDD VDD GND sky130_ef_sc_hd__decap_12
Xinput1 input1/A GND GND VDD VDD net1 sky130_fd_sc_hd__buf_2
XPHY_EDGE_ROW_9_Right_9 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_0_11_53 GND GND VDD VDD sky130_fd_sc_hd__decap_3
Xinput2 reset GND GND VDD VDD net2 sky130_fd_sc_hd__clkbuf_4
Xinput3 input3/A GND GND VDD VDD net3 sky130_fd_sc_hd__clkbuf_2
XPHY_EDGE_ROW_7_Left_19 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_0_Right_0 GND GND VDD VDD sky130_fd_sc_hd__decap_3
Xinput4 input4/A GND GND VDD VDD net4 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_5_52 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_10_Left_22 GND GND VDD VDD sky130_fd_sc_hd__decap_3
X_76_ net13 GND GND VDD VDD net14 sky130_fd_sc_hd__clkbuf_1
Xinput5 input5/A GND GND VDD VDD net5 sky130_fd_sc_hd__dlymetal6s2s_1
X_59_ _12_ net5 net10 GND GND VDD VDD _28_ sky130_fd_sc_hd__o21a_1
X_58_ _08_ _09_ net12 GND GND VDD VDD _27_ sky130_fd_sc_hd__nor3b_1
X_75_ clknet_1_1__leaf_clk net16 net2 GND GND VDD VDD net13 sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_4_Right_4 GND GND VDD VDD sky130_fd_sc_hd__decap_3
X_74_ clknet_1_1__leaf_clk _06_ net2 GND GND VDD VDD net12 sky130_fd_sc_hd__dfrtp_1
X_57_ _11_ _24_ _25_ _26_ GND GND VDD VDD _04_ sky130_fd_sc_hd__o31a_1
X_73_ clknet_1_1__leaf_clk _05_ net2 GND GND VDD VDD net11 sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_2_Left_14 GND GND VDD VDD sky130_fd_sc_hd__decap_3
X_56_ net3 net1 net10 GND GND VDD VDD _26_ sky130_fd_sc_hd__or3_1
Xclkbuf_1_0__f_clk clknet_0_clk GND GND VDD VDD clknet_1_0__leaf_clk sky130_fd_sc_hd__clkbuf_16
X_39_ _12_ net4 GND GND VDD VDD _13_ sky130_fd_sc_hd__and2_1
X_72_ clknet_1_1__leaf_clk _04_ net2 GND GND VDD VDD net10 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_5_57 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_10_Right_10 GND GND VDD VDD sky130_fd_sc_hd__decap_3
X_55_ _12_ net5 net9 GND GND VDD VDD _25_ sky130_fd_sc_hd__o21a_1
X_38_ net3 GND GND VDD VDD _12_ sky130_fd_sc_hd__buf_2
Xhold1 net12 GND GND VDD VDD net15 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_8_Right_8 GND GND VDD VDD sky130_fd_sc_hd__decap_3
X_71_ clknet_1_0__leaf_clk _03_ net2 GND GND VDD VDD net9 sky130_fd_sc_hd__dfrtp_1
X_54_ _08_ _09_ net11 GND GND VDD VDD _24_ sky130_fd_sc_hd__nor3b_1
X_37_ net3 net1 GND GND VDD VDD _11_ sky130_fd_sc_hd__nor2_2
Xhold2 _07_ GND GND VDD VDD net16 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_8_25 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_0_11_29 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_70_ clknet_1_0__leaf_clk _02_ net2 GND GND VDD VDD net8 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_5_37 GND GND VDD VDD sky130_fd_sc_hd__decap_8
X_53_ _11_ _21_ _22_ _23_ GND GND VDD VDD _03_ sky130_fd_sc_hd__o31a_1
XPHY_EDGE_ROW_6_Left_18 GND GND VDD VDD sky130_fd_sc_hd__decap_3
X_36_ _08_ _09_ net7 GND GND VDD VDD _10_ sky130_fd_sc_hd__nor3b_1
XPHY_EDGE_ROW_9_Left_21 GND GND VDD VDD sky130_fd_sc_hd__decap_3
Xhold3 net8 GND GND VDD VDD net17 sky130_fd_sc_hd__dlygate4sd3_1
X_52_ _12_ net1 net9 GND GND VDD VDD _23_ sky130_fd_sc_hd__or3_1
X_35_ net5 GND GND VDD VDD _09_ sky130_fd_sc_hd__buf_2
Xhold4 net12 GND GND VDD VDD net18 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_10_9 GND GND VDD VDD sky130_fd_sc_hd__decap_8
X_51_ _12_ net5 net8 GND GND VDD VDD _22_ sky130_fd_sc_hd__o21a_1
XFILLER_0_2_29 GND GND VDD VDD sky130_fd_sc_hd__decap_4
X_34_ net3 GND GND VDD VDD _08_ sky130_fd_sc_hd__buf_2
XFILLER_0_5_18 GND GND VDD VDD sky130_fd_sc_hd__decap_8
XFILLER_0_6_61 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_0_6_3 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_50_ _08_ _09_ net10 GND GND VDD VDD _21_ sky130_fd_sc_hd__nor3b_1
Xclkbuf_1_1__f_clk clknet_0_clk GND GND VDD VDD clknet_1_1__leaf_clk sky130_fd_sc_hd__clkbuf_16
XPHY_EDGE_ROW_3_Right_3 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_0_3_52 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_1_Left_13 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_0_4_3 GND GND VDD VDD sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_7_Right_7 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_0_0_34 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_5_Left_17 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_0_0_46 GND GND VDD VDD sky130_fd_sc_hd__decap_8
XFILLER_0_0_57 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_8_Left_20 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_0_2_3 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_0_0_15 GND VDD VDD GND sky130_ef_sc_hd__decap_12
X_69_ clknet_1_0__leaf_clk _01_ net2 GND GND VDD VDD net7 sky130_fd_sc_hd__dfrtp_1
X_68_ clknet_1_0__leaf_clk _00_ net2 GND GND VDD VDD net6 sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_2_Right_2 GND GND VDD VDD sky130_fd_sc_hd__decap_3
X_67_ _08_ net1 net13 _33_ net15 GND GND VDD VDD _07_ sky130_fd_sc_hd__o32a_1
XFILLER_0_0_3 GND VDD VDD GND sky130_ef_sc_hd__decap_12
XFILLER_0_6_49 GND VDD VDD GND sky130_ef_sc_hd__decap_12
Xoutput6 net6 GND GND VDD VDD data_out[0] sky130_fd_sc_hd__clkbuf_4
C0 _08_ VDD 2.09f
C1 VDD net1 5.95f
C2 net9 VDD 2.27f
C3 VDD clknet_1_0__leaf_clk 2.53f
C4 net2 VDD 2.2f
C5 clknet_1_1__leaf_clk VDD 2.8f
C6 _08_ _09_ 2.33f
C7 _09_ VDD 2.97f
C8 _12_ net1 2.74f
C9 net6 VDD 2.06f
C10 VDD _12_ 2.83f
C11 net2 GND 5.94f
C12 net10 GND 3.07f
C13 net8 GND 2.48f
C14 _12_ GND 3.92f
C15 net1 GND 3.49f
C16 VDD GND 0.13p
C17 clknet_0_clk GND 2.69f
C18 _11_ GND 3.4f
C19 clkbuf_0_clk/A GND 3.74f
C20 _08_ GND 2.76f
C21 net3 GND 3.25f
C22 net7 GND 3.41f
.ends

.subckt reconfigurable_CP
XCP2_5_stage_0 CP2_5_stage_0/charge_pump_reverse_1/nmos_dnw3_0/vs CP1_5_stage_0/charge_pump1_0/clk_in
+ VSUBS CP2_5_stage_0/charge_pump_reverse_1/clock_0/clk_in CP2_5_stage_1/charge_pump_0/nmos_dnw3_0/vin
+ CP2_5_stage_0/charge_pump_reverse_0/nmos_dnw3_0/vin CP1_5_stage_0/charge_pump1_2/vdd
+ scanchain_0/data_out[1] CP2_5_stage_0/charge_pump_0/nmos_dnw3_0/vin scanchain_0/data_out[6]
+ CP2_5_stage_0/charge_pump_0/nmos_dnw3_0/vs VSUBS scanchain_0/data_out[2] scanchain_0/data_out[7]
+ CP2_5_stage_0/charge_pump_2/nmos_dnw3_0/vs scanchain_0/data_out[4] CP2_5_stage_0/charge_pump_1/nmos_dnw3_0/vs
+ CP2_5_stage_0/charge_pump_reverse_0/nmos_dnw3_0/vs scanchain_0/data_out[3] CP1_5_stage_0/charge_pump1_0/clk_in
+ CP2_5_stage_0/charge_pump_0/clock_0/clk_in CP2_5_stage_0/charge_pump_reverse_1/clock_0/clk_in
+ scanchain_0/data_out[0] scanchain_0/data_out[5] VSUBS CP2_5_stage
XCP2_5_stage_1 CP2_5_stage_1/charge_pump_reverse_1/nmos_dnw3_0/vs CP2_5_stage_1/m1_94493_n2143#
+ CP2_5_stage_1/charge_pump_reverse_1/nmos_dnw3_0/out2 CP2_5_stage_1/m1_71529_n2069#
+ CP2_5_stage_1/charge_pump_2/m1_12174_n760# CP2_5_stage_1/charge_pump_reverse_0/nmos_dnw3_0/vin
+ CP1_5_stage_0/charge_pump1_2/vdd scanchain_0/data_out[6] CP2_5_stage_1/charge_pump_0/nmos_dnw3_0/vin
+ scanchain_0/data_out[1] CP2_5_stage_1/charge_pump_0/nmos_dnw3_0/vs CP2_5_stage_1/charge_pump_reverse_1/clock_0/clk
+ scanchain_0/data_out[5] scanchain_0/data_out[0] CP2_5_stage_1/charge_pump_2/nmos_dnw3_0/vs
+ scanchain_0/data_out[3] CP2_5_stage_1/charge_pump_1/nmos_dnw3_0/vs CP2_5_stage_1/charge_pump_reverse_0/nmos_dnw3_0/vs
+ scanchain_0/data_out[4] CP2_5_stage_1/charge_pump_2/clock_0/clk_in CP1_5_stage_0/charge_pump1_0/clk_in
+ CP2_5_stage_1/charge_pump_reverse_1/clock_0/clk_in scanchain_0/data_out[7] scanchain_0/data_out[2]
+ VSUBS CP2_5_stage
XCP1_5_stage_0 CP1_5_stage_0/charge_pump1_2/vdd scanchain_0/data_out[7] scanchain_0/data_out[0]
+ scanchain_0/data_out[1] CP2_5_stage_0/charge_pump_0/nmos_dnw3_0/vin scanchain_0/data_out[2]
+ CP1_5_stage_0/charge_pump1_reverse_0/nmos_dnw3_0/vs scanchain_0/data_out[3] CP1_5_stage_0/charge_pump1_1/nmos_dnw3_0/vs
+ CP1_5_stage_0/charge_pump1_0/clk_in scanchain_0/data_out[4] scanchain_0/data_out[5]
+ CP1_5_stage_0/charge_pump1_0/nmos_dnw3_0/vs scanchain_0/data_out[6] CP1_5_stage_0/charge_pump1_reverse_1/nmos_dnw3_0/vs
+ CP1_5_stage_0/charge_pump1_2/nmos_dnw3_0/vs VSUBS CP1_5_stage
Xscanchain_0 scanchain_0/VDD scanchain_0/data_out[0] scanchain_0/data_out[1] scanchain_0/data_out[2]
+ scanchain_0/data_out[3] scanchain_0/data_out[4] scanchain_0/data_out[5] scanchain_0/data_out[6]
+ scanchain_0/data_out[7] scanchain_0/scan_out VSUBS scanchain
C0 scanchain_0/data_out[1] scanchain_0/data_out[6] 2.69f
C1 scanchain_0/data_out[1] scanchain_0/data_out[0] 13.4f
C2 scanchain_0/data_out[1] scanchain_0/data_out[2] 8.23f
C3 VSUBS scanchain_0/data_out[7] 2.45f
C4 scanchain_0/data_out[2] scanchain_0/data_out[3] 9.12f
C5 scanchain_0/data_out[3] scanchain_0/data_out[4] 10.5f
C6 scanchain_0/data_out[6] scanchain_0/data_out[7] 5.47f
C7 CP1_5_stage_0/charge_pump1_2/vdd CP1_5_stage_0/charge_pump1_0/clk_in 3.04f
C8 scanchain_0/data_out[1] CP1_5_stage_0/charge_pump1_0/clk_in 2.29f
C9 scanchain_0/data_out[6] VSUBS 2.01f
C10 scanchain_0/data_out[7] scanchain_0/data_out[0] 3.24f
C11 VSUBS scanchain_0/data_out[0] 2.38f
C12 scanchain_0/data_out[5] scanchain_0/data_out[6] 8.2f
C13 CP1_5_stage_0/charge_pump1_2/vdd VSUBS 7.26f
C14 scanchain_0/data_out[5] scanchain_0/data_out[4] 9.18f
C15 scanchain_0/data_out[2] scanchain_0/data_out[6] 2.24f
C16 scanchain_0/net2 0 2.35f
C17 scanchain_0/VDD 0 88.6f
C18 scanchain_0/clkbuf_0_clk/A 0 2.59f
C19 CP1_5_stage_0/charge_pump1_reverse_1/input1 0 22.9f
C20 CP1_5_stage_0/charge_pump1_reverse_1/input2 0 22.4f
C21 CP1_5_stage_0/charge_pump1_reverse_1/capacitors_1_12/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C22 CP1_5_stage_0/charge_pump1_reverse_1/capacitors_1_12/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C23 CP1_5_stage_0/charge_pump1_reverse_1/capacitors_1_12/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 0 2.66f
C24 CP1_5_stage_0/charge_pump1_reverse_1/capacitors_1_13/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C25 CP1_5_stage_0/charge_pump1_reverse_1/capacitors_1_13/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C26 CP1_5_stage_0/charge_pump1_reverse_1/capacitors_1_13/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 0 2.66f
C27 CP1_5_stage_0/charge_pump1_reverse_1/capacitors_1_11/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C28 CP1_5_stage_0/charge_pump1_reverse_1/capacitors_1_11/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C29 CP1_5_stage_0/charge_pump1_reverse_1/capacitors_1_11/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 0 2.66f
C30 CP1_5_stage_0/charge_pump1_reverse_1/capacitors_1_10/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C31 CP1_5_stage_0/charge_pump1_reverse_1/capacitors_1_10/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C32 CP1_5_stage_0/charge_pump1_reverse_1/capacitors_1_10/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 0 2.66f
C33 CP1_5_stage_0/charge_pump1_reverse_1/m1_4341_n519# 0 3.86f
C34 CP1_5_stage_0/charge_pump1_reverse_1/m1_12659_300# 0 2.73f
C35 CP1_5_stage_0/charge_pump1_2/nmos_dnw3_0/vs 0 15.1f
C36 CP1_5_stage_0/charge_pump1_reverse_1/capacitors_1_9/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C37 CP1_5_stage_0/charge_pump1_reverse_1/capacitors_1_9/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C38 CP1_5_stage_0/charge_pump1_reverse_1/capacitors_1_9/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 0 2.66f
C39 CP1_5_stage_0/charge_pump1_reverse_1/capacitors_1_8/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C40 CP1_5_stage_0/charge_pump1_reverse_1/capacitors_1_8/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C41 CP1_5_stage_0/charge_pump1_reverse_1/capacitors_1_8/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 0 2.66f
C42 CP1_5_stage_0/charge_pump1_reverse_1/capacitors_1_7/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C43 CP1_5_stage_0/charge_pump1_reverse_1/capacitors_1_7/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C44 CP1_5_stage_0/charge_pump1_reverse_1/capacitors_1_7/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 0 2.66f
C45 CP1_5_stage_0/charge_pump1_reverse_1/capacitors_1_6/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C46 CP1_5_stage_0/charge_pump1_reverse_1/capacitors_1_6/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C47 CP1_5_stage_0/charge_pump1_reverse_1/capacitors_1_6/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 0 2.66f
C48 CP1_5_stage_0/charge_pump1_reverse_1/capacitors_1_5/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C49 CP1_5_stage_0/charge_pump1_reverse_1/capacitors_1_5/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C50 CP1_5_stage_0/charge_pump1_reverse_1/capacitors_1_5/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 0 2.66f
C51 CP1_5_stage_0/charge_pump1_reverse_1/capacitors_1_4/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C52 CP1_5_stage_0/charge_pump1_reverse_1/capacitors_1_4/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C53 CP1_5_stage_0/charge_pump1_reverse_1/capacitors_1_4/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 0 2.66f
C54 CP1_5_stage_0/charge_pump1_reverse_1/capacitors_1_3/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C55 CP1_5_stage_0/charge_pump1_reverse_1/capacitors_1_3/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C56 CP1_5_stage_0/charge_pump1_reverse_1/capacitors_1_3/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 0 2.66f
C57 CP1_5_stage_0/charge_pump1_reverse_1/capacitors_1_2/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C58 CP1_5_stage_0/charge_pump1_reverse_1/capacitors_1_2/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C59 CP1_5_stage_0/charge_pump1_reverse_1/capacitors_1_2/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 0 2.66f
C60 CP1_5_stage_0/charge_pump1_reverse_1/capacitors_1_1/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C61 CP1_5_stage_0/charge_pump1_reverse_1/capacitors_1_1/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C62 CP1_5_stage_0/charge_pump1_reverse_1/capacitors_1_1/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 0 2.66f
C63 CP1_5_stage_0/charge_pump1_reverse_1/capacitors_1_0/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C64 CP1_5_stage_0/charge_pump1_reverse_1/capacitors_1_0/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C65 CP1_5_stage_0/charge_pump1_reverse_1/capacitors_1_0/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 0 2.66f
C66 CP1_5_stage_0/charge_pump1_reverse_1/capacitor_8_1/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C67 CP1_5_stage_0/charge_pump1_reverse_1/clock_1/clk 0 88.1f
C68 CP1_5_stage_0/charge_pump1_reverse_1/capacitor_8_1/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C69 CP1_5_stage_0/charge_pump1_reverse_1/capacitor_8_1/capacitor_7_0/buffer_and_gate_0/in1 0 2.66f
C70 CP1_5_stage_0/charge_pump1_reverse_1/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C71 CP1_5_stage_0/charge_pump1_reverse_1/clock_1/clkb 0 96.8f
C72 CP1_5_stage_0/charge_pump1_reverse_1/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C73 CP1_5_stage_0/charge_pump1_reverse_1/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 0 2.66f
C74 CP1_5_stage_0/charge_pump1_reverse_1/clock_1/a_2432_n962# 0 8.68f **FLOATING
C75 CP1_5_stage_0/charge_pump1_reverse_1/clock_1/a_2020_n482# 0 2.57f **FLOATING
C76 CP1_5_stage_0/charge_pump1_reverse_1/clock_1/a_344_102# 0 2.81f
C77 CP1_5_stage_0/charge_pump1_reverse_1/clock_1/a_2402_572# 0 2.17f
C78 CP1_5_stage_0/charge_pump1_reverse_1/clock_1/a_344_n986# 0 2.38f
C79 CP1_5_stage_0/charge_pump1_reverse_1/clock_1/clk_in 0 14.7f
C80 CP1_5_stage_0/charge_pump1_reverse_1/clock_1/a_3246_118# 0 6.83f
C81 CP1_5_stage_0/charge_pump1_reverse_1/nmos_dnw3_0/clkb 0 2.01f
C82 CP1_5_stage_0/charge_pump1_reverse_0/input1 0 22.9f
C83 CP1_5_stage_0/charge_pump1_reverse_0/input2 0 22.4f
C84 CP1_5_stage_0/charge_pump1_reverse_0/capacitors_1_12/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C85 CP1_5_stage_0/charge_pump1_reverse_0/capacitors_1_12/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C86 CP1_5_stage_0/charge_pump1_reverse_0/capacitors_1_12/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 0 2.66f
C87 CP1_5_stage_0/charge_pump1_reverse_0/capacitors_1_13/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C88 CP1_5_stage_0/charge_pump1_reverse_0/capacitors_1_13/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C89 CP1_5_stage_0/charge_pump1_reverse_0/capacitors_1_13/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 0 2.66f
C90 CP1_5_stage_0/charge_pump1_reverse_0/capacitors_1_11/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C91 CP1_5_stage_0/charge_pump1_reverse_0/capacitors_1_11/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C92 CP1_5_stage_0/charge_pump1_reverse_0/capacitors_1_11/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 0 2.66f
C93 CP1_5_stage_0/charge_pump1_reverse_0/capacitors_1_10/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C94 CP1_5_stage_0/charge_pump1_reverse_0/capacitors_1_10/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C95 CP1_5_stage_0/charge_pump1_reverse_0/capacitors_1_10/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 0 2.66f
C96 CP1_5_stage_0/charge_pump1_reverse_0/m1_4341_n519# 0 3.86f
C97 CP1_5_stage_0/charge_pump1_reverse_0/m1_12659_300# 0 2.73f
C98 CP1_5_stage_0/charge_pump1_1/nmos_dnw3_0/vs 0 15.1f
C99 CP1_5_stage_0/charge_pump1_reverse_0/capacitors_1_9/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C100 CP1_5_stage_0/charge_pump1_reverse_0/capacitors_1_9/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C101 CP1_5_stage_0/charge_pump1_reverse_0/capacitors_1_9/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 0 2.66f
C102 CP1_5_stage_0/charge_pump1_reverse_0/capacitors_1_8/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C103 CP1_5_stage_0/charge_pump1_reverse_0/capacitors_1_8/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C104 CP1_5_stage_0/charge_pump1_reverse_0/capacitors_1_8/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 0 2.66f
C105 CP1_5_stage_0/charge_pump1_reverse_0/capacitors_1_7/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C106 CP1_5_stage_0/charge_pump1_reverse_0/capacitors_1_7/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C107 CP1_5_stage_0/charge_pump1_reverse_0/capacitors_1_7/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 0 2.66f
C108 CP1_5_stage_0/charge_pump1_reverse_0/capacitors_1_6/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C109 CP1_5_stage_0/charge_pump1_reverse_0/capacitors_1_6/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C110 CP1_5_stage_0/charge_pump1_reverse_0/capacitors_1_6/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 0 2.66f
C111 CP1_5_stage_0/charge_pump1_reverse_0/capacitors_1_5/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C112 CP1_5_stage_0/charge_pump1_reverse_0/capacitors_1_5/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C113 CP1_5_stage_0/charge_pump1_reverse_0/capacitors_1_5/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 0 2.66f
C114 CP1_5_stage_0/charge_pump1_reverse_0/capacitors_1_4/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C115 CP1_5_stage_0/charge_pump1_reverse_0/capacitors_1_4/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C116 CP1_5_stage_0/charge_pump1_reverse_0/capacitors_1_4/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 0 2.66f
C117 CP1_5_stage_0/charge_pump1_reverse_0/capacitors_1_3/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C118 CP1_5_stage_0/charge_pump1_reverse_0/capacitors_1_3/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C119 CP1_5_stage_0/charge_pump1_reverse_0/capacitors_1_3/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 0 2.66f
C120 CP1_5_stage_0/charge_pump1_reverse_0/capacitors_1_2/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C121 CP1_5_stage_0/charge_pump1_reverse_0/capacitors_1_2/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C122 CP1_5_stage_0/charge_pump1_reverse_0/capacitors_1_2/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 0 2.66f
C123 CP1_5_stage_0/charge_pump1_reverse_0/capacitors_1_1/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C124 CP1_5_stage_0/charge_pump1_reverse_0/capacitors_1_1/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C125 CP1_5_stage_0/charge_pump1_reverse_0/capacitors_1_1/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 0 2.66f
C126 CP1_5_stage_0/charge_pump1_reverse_0/capacitors_1_0/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C127 CP1_5_stage_0/charge_pump1_reverse_0/capacitors_1_0/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C128 CP1_5_stage_0/charge_pump1_reverse_0/capacitors_1_0/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 0 2.66f
C129 CP1_5_stage_0/charge_pump1_reverse_0/capacitor_8_1/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C130 CP1_5_stage_0/charge_pump1_reverse_0/clock_1/clk 0 88.1f
C131 CP1_5_stage_0/charge_pump1_reverse_0/capacitor_8_1/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C132 CP1_5_stage_0/charge_pump1_reverse_0/capacitor_8_1/capacitor_7_0/buffer_and_gate_0/in1 0 2.66f
C133 CP1_5_stage_0/charge_pump1_reverse_0/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C134 CP1_5_stage_0/charge_pump1_reverse_0/clock_1/clkb 0 96.8f
C135 CP1_5_stage_0/charge_pump1_reverse_0/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C136 CP1_5_stage_0/charge_pump1_reverse_0/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 0 2.66f
C137 CP1_5_stage_0/charge_pump1_reverse_0/clock_1/a_2432_n962# 0 8.68f **FLOATING
C138 CP1_5_stage_0/charge_pump1_reverse_0/clock_1/a_2020_n482# 0 2.57f **FLOATING
C139 CP1_5_stage_0/charge_pump1_reverse_0/clock_1/a_344_102# 0 2.81f
C140 CP1_5_stage_0/charge_pump1_reverse_0/clock_1/a_2402_572# 0 2.17f
C141 CP1_5_stage_0/charge_pump1_reverse_0/clock_1/a_344_n986# 0 2.38f
C142 CP1_5_stage_0/charge_pump1_reverse_0/clock_1/clk_in 0 12.2f
C143 CP1_5_stage_0/charge_pump1_reverse_0/clock_1/a_3246_118# 0 6.83f
C144 CP1_5_stage_0/charge_pump1_reverse_0/nmos_dnw3_0/clkb 0 2.01f
C145 CP1_5_stage_0/charge_pump1_2/input1 0 22.5f
C146 CP1_5_stage_0/charge_pump1_2/input2 0 22.2f
C147 CP1_5_stage_0/charge_pump1_2/capacitors_1_12/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C148 CP1_5_stage_0/charge_pump1_2/capacitors_1_12/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C149 CP1_5_stage_0/charge_pump1_2/capacitors_1_12/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 0 2.66f
C150 CP1_5_stage_0/charge_pump1_2/capacitors_1_13/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C151 CP1_5_stage_0/charge_pump1_2/capacitors_1_13/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C152 CP1_5_stage_0/charge_pump1_2/capacitors_1_13/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 0 2.66f
C153 CP1_5_stage_0/charge_pump1_2/capacitors_1_11/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C154 CP1_5_stage_0/charge_pump1_2/capacitors_1_11/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C155 CP1_5_stage_0/charge_pump1_2/capacitors_1_11/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 0 2.66f
C156 CP1_5_stage_0/charge_pump1_2/capacitors_1_10/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C157 CP1_5_stage_0/charge_pump1_2/capacitors_1_10/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C158 CP1_5_stage_0/charge_pump1_2/capacitors_1_10/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 0 2.66f
C159 CP1_5_stage_0/charge_pump1_2/m1_4341_n519# 0 3.77f
C160 CP1_5_stage_0/charge_pump1_2/m1_12659_300# 0 2.54f
C161 CP2_5_stage_0/charge_pump_0/nmos_dnw3_0/vin 0 5.86f
C162 CP1_5_stage_0/charge_pump1_2/capacitors_1_9/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C163 CP1_5_stage_0/charge_pump1_2/capacitors_1_9/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C164 CP1_5_stage_0/charge_pump1_2/capacitors_1_9/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 0 2.66f
C165 CP1_5_stage_0/charge_pump1_2/capacitors_1_8/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C166 CP1_5_stage_0/charge_pump1_2/capacitors_1_8/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C167 CP1_5_stage_0/charge_pump1_2/capacitors_1_8/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 0 2.66f
C168 CP1_5_stage_0/charge_pump1_2/capacitors_1_7/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C169 CP1_5_stage_0/charge_pump1_2/capacitors_1_7/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C170 CP1_5_stage_0/charge_pump1_2/capacitors_1_7/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 0 2.66f
C171 CP1_5_stage_0/charge_pump1_2/capacitors_1_6/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C172 CP1_5_stage_0/charge_pump1_2/capacitors_1_6/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C173 CP1_5_stage_0/charge_pump1_2/capacitors_1_6/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 0 2.66f
C174 CP1_5_stage_0/charge_pump1_2/capacitors_1_5/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C175 CP1_5_stage_0/charge_pump1_2/capacitors_1_5/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C176 CP1_5_stage_0/charge_pump1_2/capacitors_1_5/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 0 2.66f
C177 CP1_5_stage_0/charge_pump1_2/capacitors_1_4/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C178 CP1_5_stage_0/charge_pump1_2/capacitors_1_4/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C179 CP1_5_stage_0/charge_pump1_2/capacitors_1_4/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 0 2.66f
C180 CP1_5_stage_0/charge_pump1_2/capacitors_1_3/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C181 CP1_5_stage_0/charge_pump1_2/capacitors_1_3/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C182 CP1_5_stage_0/charge_pump1_2/capacitors_1_3/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 0 2.66f
C183 CP1_5_stage_0/charge_pump1_2/capacitors_1_2/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C184 CP1_5_stage_0/charge_pump1_2/capacitors_1_2/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C185 CP1_5_stage_0/charge_pump1_2/capacitors_1_2/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 0 2.66f
C186 CP1_5_stage_0/charge_pump1_2/capacitors_1_1/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C187 CP1_5_stage_0/charge_pump1_2/capacitors_1_1/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C188 CP1_5_stage_0/charge_pump1_2/capacitors_1_1/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 0 2.66f
C189 CP1_5_stage_0/charge_pump1_2/capacitors_1_0/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C190 CP1_5_stage_0/charge_pump1_2/capacitors_1_0/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C191 CP1_5_stage_0/charge_pump1_2/capacitors_1_0/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 0 2.66f
C192 CP1_5_stage_0/charge_pump1_2/capacitor_8_1/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C193 CP1_5_stage_0/charge_pump1_2/clock_0/clkb 0 86.1f
C194 CP1_5_stage_0/charge_pump1_2/capacitor_8_1/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C195 CP1_5_stage_0/charge_pump1_2/capacitor_8_1/capacitor_7_0/buffer_and_gate_0/in1 0 2.66f
C196 CP1_5_stage_0/charge_pump1_2/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C197 CP1_5_stage_0/charge_pump1_2/clock_0/clk 0 85.5f
C198 CP1_5_stage_0/charge_pump1_2/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C199 CP1_5_stage_0/charge_pump1_2/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 0 2.66f
C200 CP1_5_stage_0/charge_pump1_2/clock_0/a_2432_n962# 0 8.68f **FLOATING
C201 CP1_5_stage_0/charge_pump1_2/clock_0/a_2020_n482# 0 2.57f **FLOATING
C202 CP1_5_stage_0/charge_pump1_2/clock_0/a_344_102# 0 2.81f
C203 CP1_5_stage_0/charge_pump1_2/clock_0/a_2402_572# 0 2.17f
C204 CP1_5_stage_0/charge_pump1_2/clock_0/a_344_n986# 0 2.38f
C205 CP1_5_stage_0/charge_pump1_2/clk_in 0 11.3f
C206 CP1_5_stage_0/charge_pump1_2/clock_0/a_3246_118# 0 6.83f
C207 CP1_5_stage_0/charge_pump1_2/nmos_dnw3_0/clkb 0 2.34f
C208 CP1_5_stage_0/charge_pump1_1/input1 0 22.5f
C209 CP1_5_stage_0/charge_pump1_1/input2 0 22.2f
C210 CP1_5_stage_0/charge_pump1_1/capacitors_1_12/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C211 CP1_5_stage_0/charge_pump1_1/capacitors_1_12/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C212 CP1_5_stage_0/charge_pump1_1/capacitors_1_12/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 0 2.66f
C213 CP1_5_stage_0/charge_pump1_1/capacitors_1_13/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C214 CP1_5_stage_0/charge_pump1_1/capacitors_1_13/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C215 CP1_5_stage_0/charge_pump1_1/capacitors_1_13/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 0 2.66f
C216 CP1_5_stage_0/charge_pump1_1/capacitors_1_11/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C217 CP1_5_stage_0/charge_pump1_1/capacitors_1_11/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C218 CP1_5_stage_0/charge_pump1_1/capacitors_1_11/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 0 2.66f
C219 CP1_5_stage_0/charge_pump1_1/capacitors_1_10/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C220 CP1_5_stage_0/charge_pump1_1/capacitors_1_10/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C221 CP1_5_stage_0/charge_pump1_1/capacitors_1_10/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 0 2.66f
C222 CP1_5_stage_0/charge_pump1_1/m1_4341_n519# 0 3.77f
C223 CP1_5_stage_0/charge_pump1_1/m1_12659_300# 0 2.54f
C224 CP1_5_stage_0/charge_pump1_reverse_1/nmos_dnw3_0/vs 0 14.5f
C225 CP1_5_stage_0/charge_pump1_1/capacitors_1_9/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C226 CP1_5_stage_0/charge_pump1_1/capacitors_1_9/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C227 CP1_5_stage_0/charge_pump1_1/capacitors_1_9/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 0 2.66f
C228 CP1_5_stage_0/charge_pump1_1/capacitors_1_8/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C229 CP1_5_stage_0/charge_pump1_1/capacitors_1_8/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C230 CP1_5_stage_0/charge_pump1_1/capacitors_1_8/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 0 2.66f
C231 CP1_5_stage_0/charge_pump1_1/capacitors_1_7/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C232 CP1_5_stage_0/charge_pump1_1/capacitors_1_7/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C233 CP1_5_stage_0/charge_pump1_1/capacitors_1_7/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 0 2.66f
C234 CP1_5_stage_0/charge_pump1_1/capacitors_1_6/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C235 CP1_5_stage_0/charge_pump1_1/capacitors_1_6/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C236 CP1_5_stage_0/charge_pump1_1/capacitors_1_6/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 0 2.66f
C237 CP1_5_stage_0/charge_pump1_1/capacitors_1_5/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C238 CP1_5_stage_0/charge_pump1_1/capacitors_1_5/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C239 CP1_5_stage_0/charge_pump1_1/capacitors_1_5/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 0 2.66f
C240 CP1_5_stage_0/charge_pump1_1/capacitors_1_4/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C241 CP1_5_stage_0/charge_pump1_1/capacitors_1_4/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C242 CP1_5_stage_0/charge_pump1_1/capacitors_1_4/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 0 2.66f
C243 CP1_5_stage_0/charge_pump1_1/capacitors_1_3/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C244 CP1_5_stage_0/charge_pump1_1/capacitors_1_3/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C245 CP1_5_stage_0/charge_pump1_1/capacitors_1_3/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 0 2.66f
C246 CP1_5_stage_0/charge_pump1_1/capacitors_1_2/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C247 CP1_5_stage_0/charge_pump1_1/capacitors_1_2/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C248 CP1_5_stage_0/charge_pump1_1/capacitors_1_2/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 0 2.66f
C249 CP1_5_stage_0/charge_pump1_1/capacitors_1_1/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C250 CP1_5_stage_0/charge_pump1_1/capacitors_1_1/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C251 CP1_5_stage_0/charge_pump1_1/capacitors_1_1/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 0 2.66f
C252 CP1_5_stage_0/charge_pump1_1/capacitors_1_0/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C253 CP1_5_stage_0/charge_pump1_1/capacitors_1_0/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C254 CP1_5_stage_0/charge_pump1_1/capacitors_1_0/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 0 2.66f
C255 CP1_5_stage_0/charge_pump1_1/capacitor_8_1/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C256 CP1_5_stage_0/charge_pump1_1/clock_0/clkb 0 86.1f
C257 CP1_5_stage_0/charge_pump1_1/capacitor_8_1/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C258 CP1_5_stage_0/charge_pump1_1/capacitor_8_1/capacitor_7_0/buffer_and_gate_0/in1 0 2.66f
C259 CP1_5_stage_0/charge_pump1_1/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C260 CP1_5_stage_0/charge_pump1_1/clock_0/clk 0 85.5f
C261 CP1_5_stage_0/charge_pump1_1/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C262 CP1_5_stage_0/charge_pump1_1/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 0 2.66f
C263 CP1_5_stage_0/charge_pump1_1/clock_0/a_2432_n962# 0 8.68f **FLOATING
C264 CP1_5_stage_0/charge_pump1_1/clock_0/a_2020_n482# 0 2.57f **FLOATING
C265 CP1_5_stage_0/charge_pump1_1/clock_0/a_344_102# 0 2.81f
C266 CP1_5_stage_0/charge_pump1_1/clock_0/a_2402_572# 0 2.17f
C267 CP1_5_stage_0/charge_pump1_1/clock_0/a_344_n986# 0 2.38f
C268 CP1_5_stage_0/charge_pump1_1/clk_in 0 18.2f
C269 CP1_5_stage_0/charge_pump1_1/clock_0/a_3246_118# 0 6.83f
C270 CP1_5_stage_0/charge_pump1_1/nmos_dnw3_0/clkb 0 2.34f
C271 CP1_5_stage_0/charge_pump1_0/input1 0 22.5f
C272 CP1_5_stage_0/charge_pump1_0/input2 0 22.2f
C273 CP1_5_stage_0/charge_pump1_0/capacitors_1_12/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C274 CP1_5_stage_0/charge_pump1_0/capacitors_1_12/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C275 CP1_5_stage_0/charge_pump1_0/capacitors_1_12/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 0 2.66f
C276 CP1_5_stage_0/charge_pump1_0/capacitors_1_13/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C277 CP1_5_stage_0/charge_pump1_0/capacitors_1_13/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C278 CP1_5_stage_0/charge_pump1_0/capacitors_1_13/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 0 2.66f
C279 CP1_5_stage_0/charge_pump1_0/capacitors_1_11/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C280 CP1_5_stage_0/charge_pump1_0/capacitors_1_11/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C281 CP1_5_stage_0/charge_pump1_0/capacitors_1_11/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 0 2.66f
C282 CP1_5_stage_0/charge_pump1_0/capacitors_1_10/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C283 CP1_5_stage_0/charge_pump1_0/capacitors_1_10/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C284 CP1_5_stage_0/charge_pump1_0/capacitors_1_10/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 0 2.66f
C285 CP1_5_stage_0/charge_pump1_0/m1_4341_n519# 0 3.77f
C286 CP1_5_stage_0/charge_pump1_0/m1_12659_300# 0 2.54f
C287 CP1_5_stage_0/charge_pump1_reverse_0/nmos_dnw3_0/vs 0 14.7f
C288 CP1_5_stage_0/charge_pump1_0/capacitors_1_9/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C289 CP1_5_stage_0/charge_pump1_0/capacitors_1_9/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C290 CP1_5_stage_0/charge_pump1_0/capacitors_1_9/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 0 2.66f
C291 CP1_5_stage_0/charge_pump1_0/capacitors_1_8/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C292 CP1_5_stage_0/charge_pump1_0/capacitors_1_8/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C293 CP1_5_stage_0/charge_pump1_0/capacitors_1_8/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 0 2.66f
C294 CP1_5_stage_0/charge_pump1_0/capacitors_1_7/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C295 CP1_5_stage_0/charge_pump1_0/capacitors_1_7/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C296 CP1_5_stage_0/charge_pump1_0/capacitors_1_7/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 0 2.66f
C297 CP1_5_stage_0/charge_pump1_0/capacitors_1_6/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C298 CP1_5_stage_0/charge_pump1_0/capacitors_1_6/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C299 CP1_5_stage_0/charge_pump1_0/capacitors_1_6/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 0 2.66f
C300 CP1_5_stage_0/charge_pump1_0/capacitors_1_5/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C301 CP1_5_stage_0/charge_pump1_0/capacitors_1_5/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C302 CP1_5_stage_0/charge_pump1_0/capacitors_1_5/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 0 2.66f
C303 CP1_5_stage_0/charge_pump1_0/capacitors_1_4/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C304 CP1_5_stage_0/charge_pump1_0/capacitors_1_4/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C305 CP1_5_stage_0/charge_pump1_0/capacitors_1_4/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 0 2.66f
C306 CP1_5_stage_0/charge_pump1_0/capacitors_1_3/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C307 CP1_5_stage_0/charge_pump1_0/capacitors_1_3/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C308 CP1_5_stage_0/charge_pump1_0/capacitors_1_3/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 0 2.66f
C309 CP1_5_stage_0/charge_pump1_0/capacitors_1_2/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C310 CP1_5_stage_0/charge_pump1_0/capacitors_1_2/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C311 CP1_5_stage_0/charge_pump1_0/capacitors_1_2/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 0 2.66f
C312 CP1_5_stage_0/charge_pump1_0/capacitors_1_1/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C313 CP1_5_stage_0/charge_pump1_0/capacitors_1_1/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C314 CP1_5_stage_0/charge_pump1_0/capacitors_1_1/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 0 2.66f
C315 CP1_5_stage_0/charge_pump1_0/capacitors_1_0/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C316 CP1_5_stage_0/charge_pump1_0/capacitors_1_0/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C317 CP1_5_stage_0/charge_pump1_0/capacitors_1_0/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 0 2.66f
C318 CP1_5_stage_0/charge_pump1_0/capacitor_8_1/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C319 CP1_5_stage_0/charge_pump1_0/clock_0/clkb 0 86.1f
C320 CP1_5_stage_0/charge_pump1_0/capacitor_8_1/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C321 CP1_5_stage_0/charge_pump1_0/capacitor_8_1/capacitor_7_0/buffer_and_gate_0/in1 0 2.66f
C322 CP1_5_stage_0/charge_pump1_0/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C323 CP1_5_stage_0/charge_pump1_0/clock_0/clk 0 85.5f
C324 CP1_5_stage_0/charge_pump1_0/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C325 CP1_5_stage_0/charge_pump1_0/capacitor_8_0/capacitor_7_0/buffer_and_gate_0/in1 0 2.66f
C326 CP1_5_stage_0/charge_pump1_0/clock_0/a_2432_n962# 0 8.68f **FLOATING
C327 CP1_5_stage_0/charge_pump1_0/clock_0/a_2020_n482# 0 2.57f **FLOATING
C328 CP1_5_stage_0/charge_pump1_0/clock_0/a_344_102# 0 2.81f
C329 CP1_5_stage_0/charge_pump1_0/clock_0/a_2402_572# 0 2.17f
C330 CP1_5_stage_0/charge_pump1_0/clock_0/a_344_n986# 0 2.38f
C331 CP1_5_stage_0/charge_pump1_0/clock_0/a_3246_118# 0 6.83f
C332 CP1_5_stage_0/charge_pump1_0/nmos_dnw3_0/clkb 0 2.34f
C333 CP1_5_stage_0/charge_pump1_0/nmos_dnw3_0/vs 0 10.4f
C334 CP2_5_stage_1/charge_pump_reverse_1/nmos_dnw3_0/vs 0 16.4f
C335 CP2_5_stage_1/charge_pump_reverse_1/sky130_fd_pr__pfet_01v8_4RPJ49_1/w_n3905_n142# 0 6.63f
C336 CP2_5_stage_1/charge_pump_reverse_1/sky130_fd_pr__pfet_01v8_4RPJ49_0/w_n3905_n142# 0 6.63f
C337 CP2_5_stage_1/charge_pump_reverse_1/clock_0/a_2432_n962# 0 8.68f **FLOATING
C338 CP2_5_stage_1/charge_pump_reverse_1/clock_0/a_2020_n482# 0 2.57f **FLOATING
C339 CP2_5_stage_1/charge_pump_reverse_1/clock_0/a_344_102# 0 2.81f
C340 CP2_5_stage_1/charge_pump_reverse_1/clock_0/a_2402_572# 0 2.17f
C341 CP2_5_stage_1/charge_pump_reverse_1/clock_0/a_344_n986# 0 2.38f
C342 CP2_5_stage_1/charge_pump_reverse_1/clock_0/a_3246_118# 0 6.83f
C343 CP2_5_stage_1/charge_pump_reverse_1/nmos_dnw3_0/clkb 0 2.23f
C344 CP2_5_stage_1/charge_pump_reverse_1/capacitors_5_0/capacitor_5_4/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C345 CP2_5_stage_1/charge_pump_reverse_1/capacitors_5_0/capacitor_5_4/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C346 CP2_5_stage_1/charge_pump_reverse_1/capacitors_5_0/capacitor_5_4/buffer_and_gate_0/in1 0 2.57f
C347 CP2_5_stage_1/charge_pump_reverse_1/capacitors_5_0/capacitor_5_3/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C348 CP2_5_stage_1/charge_pump_reverse_1/capacitors_5_0/capacitor_5_3/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C349 CP2_5_stage_1/charge_pump_reverse_1/capacitors_5_0/capacitor_5_3/buffer_and_gate_0/in1 0 2.57f
C350 CP2_5_stage_1/charge_pump_reverse_1/capacitors_5_0/capacitor_5_2/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C351 CP2_5_stage_1/charge_pump_reverse_1/capacitors_5_0/capacitor_5_2/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C352 CP2_5_stage_1/charge_pump_reverse_1/capacitors_5_0/capacitor_5_2/buffer_and_gate_0/in1 0 2.57f
C353 CP2_5_stage_1/charge_pump_reverse_1/capacitors_5_0/capacitor_5_1/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C354 CP2_5_stage_1/charge_pump_reverse_1/capacitors_5_0/capacitor_5_1/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C355 CP2_5_stage_1/charge_pump_reverse_1/capacitors_5_0/capacitor_5_1/buffer_and_gate_0/in1 0 2.57f
C356 CP2_5_stage_1/charge_pump_reverse_1/capacitors_5_0/capacitor_5_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C357 CP2_5_stage_1/charge_pump_reverse_1/capacitors_5_0/capacitor_5_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C358 CP2_5_stage_1/charge_pump_reverse_1/capacitors_5_0/capacitor_5_0/buffer_and_gate_0/in1 0 2.57f
C359 CP2_5_stage_1/charge_pump_reverse_1/nmos_dnw3_0/out1 0 15.1f
C360 CP2_5_stage_1/charge_pump_reverse_1/capacitors_5_0/capacitor_5_7/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C361 CP2_5_stage_1/charge_pump_reverse_1/clock_0/clkb 0 86.4f
C362 CP2_5_stage_1/charge_pump_reverse_1/capacitors_5_0/capacitor_5_7/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C363 CP2_5_stage_1/charge_pump_reverse_1/capacitors_5_0/capacitor_5_7/buffer_and_gate_0/in1 0 2.57f
C364 CP2_5_stage_1/charge_pump_reverse_1/capacitors_5_0/capacitor_5_6/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C365 CP2_5_stage_1/charge_pump_reverse_1/capacitors_5_0/capacitor_5_6/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C366 CP2_5_stage_1/charge_pump_reverse_1/capacitors_5_0/capacitor_5_6/buffer_and_gate_0/in1 0 2.57f
C367 CP2_5_stage_1/charge_pump_reverse_1/capacitors_5_0/capacitor_5_5/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C368 CP2_5_stage_1/charge_pump_reverse_1/capacitors_5_0/capacitor_5_5/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C369 CP2_5_stage_1/charge_pump_reverse_1/capacitors_5_0/capacitor_5_5/buffer_and_gate_0/in1 0 2.57f
C370 CP2_5_stage_1/charge_pump_reverse_1/capacitors_5_1/capacitor_5_4/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C371 CP2_5_stage_1/charge_pump_reverse_1/capacitors_5_1/capacitor_5_4/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C372 CP2_5_stage_1/charge_pump_reverse_1/capacitors_5_1/capacitor_5_4/buffer_and_gate_0/in1 0 2.57f
C373 CP2_5_stage_1/charge_pump_reverse_1/capacitors_5_1/capacitor_5_3/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C374 CP2_5_stage_1/charge_pump_reverse_1/capacitors_5_1/capacitor_5_3/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C375 CP2_5_stage_1/charge_pump_reverse_1/capacitors_5_1/capacitor_5_3/buffer_and_gate_0/in1 0 2.57f
C376 CP2_5_stage_1/charge_pump_reverse_1/capacitors_5_1/capacitor_5_2/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C377 CP2_5_stage_1/charge_pump_reverse_1/capacitors_5_1/capacitor_5_2/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C378 CP2_5_stage_1/charge_pump_reverse_1/capacitors_5_1/capacitor_5_2/buffer_and_gate_0/in1 0 2.57f
C379 CP2_5_stage_1/charge_pump_reverse_1/capacitors_5_1/capacitor_5_1/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C380 CP2_5_stage_1/charge_pump_reverse_1/capacitors_5_1/capacitor_5_1/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C381 CP2_5_stage_1/charge_pump_reverse_1/capacitors_5_1/capacitor_5_1/buffer_and_gate_0/in1 0 2.57f
C382 CP2_5_stage_1/charge_pump_reverse_1/capacitors_5_1/capacitor_5_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C383 CP2_5_stage_1/charge_pump_reverse_1/capacitors_5_1/capacitor_5_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C384 CP2_5_stage_1/charge_pump_reverse_1/capacitors_5_1/capacitor_5_0/buffer_and_gate_0/in1 0 2.57f
C385 CP2_5_stage_1/charge_pump_reverse_1/nmos_dnw3_0/out2 0 14.9f
C386 CP2_5_stage_1/charge_pump_reverse_1/capacitors_5_1/capacitor_5_7/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C387 CP2_5_stage_1/charge_pump_reverse_1/clock_0/clk 0 80f
C388 CP2_5_stage_1/charge_pump_reverse_1/capacitors_5_1/capacitor_5_7/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C389 CP2_5_stage_1/charge_pump_reverse_1/capacitors_5_1/capacitor_5_7/buffer_and_gate_0/in1 0 2.57f
C390 CP2_5_stage_1/charge_pump_reverse_1/capacitors_5_1/capacitor_5_6/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C391 CP2_5_stage_1/charge_pump_reverse_1/capacitors_5_1/capacitor_5_6/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C392 CP2_5_stage_1/charge_pump_reverse_1/capacitors_5_1/capacitor_5_6/buffer_and_gate_0/in1 0 2.57f
C393 CP2_5_stage_1/charge_pump_reverse_1/capacitors_5_1/capacitor_5_5/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C394 CP2_5_stage_1/charge_pump_reverse_1/capacitors_5_1/capacitor_5_5/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C395 CP2_5_stage_1/charge_pump_reverse_1/capacitors_5_1/capacitor_5_5/buffer_and_gate_0/in1 0 2.57f
C396 CP2_5_stage_1/charge_pump_reverse_1/nmos_dnw3_0/clk 0 2.43f
C397 CP2_5_stage_1/charge_pump_reverse_0/nmos_dnw3_0/vs 0 16.4f
C398 CP2_5_stage_1/charge_pump_reverse_0/sky130_fd_pr__pfet_01v8_4RPJ49_1/w_n3905_n142# 0 6.63f
C399 CP2_5_stage_1/charge_pump_reverse_0/sky130_fd_pr__pfet_01v8_4RPJ49_0/w_n3905_n142# 0 6.63f
C400 CP2_5_stage_1/charge_pump_reverse_0/clock_0/a_2432_n962# 0 8.68f **FLOATING
C401 CP2_5_stage_1/charge_pump_reverse_0/clock_0/a_2020_n482# 0 2.57f **FLOATING
C402 CP2_5_stage_1/charge_pump_reverse_0/clock_0/a_344_102# 0 2.81f
C403 CP2_5_stage_1/charge_pump_reverse_0/clock_0/a_2402_572# 0 2.17f
C404 CP2_5_stage_1/charge_pump_reverse_0/clock_0/a_344_n986# 0 2.38f
C405 CP2_5_stage_1/charge_pump_reverse_0/clock_0/a_3246_118# 0 6.83f
C406 CP2_5_stage_1/charge_pump_reverse_0/nmos_dnw3_0/clkb 0 2.23f
C407 CP2_5_stage_1/charge_pump_reverse_0/capacitors_5_0/capacitor_5_4/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C408 CP2_5_stage_1/charge_pump_reverse_0/capacitors_5_0/capacitor_5_4/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C409 CP2_5_stage_1/charge_pump_reverse_0/capacitors_5_0/capacitor_5_4/buffer_and_gate_0/in1 0 2.57f
C410 CP2_5_stage_1/charge_pump_reverse_0/capacitors_5_0/capacitor_5_3/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C411 CP2_5_stage_1/charge_pump_reverse_0/capacitors_5_0/capacitor_5_3/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C412 CP2_5_stage_1/charge_pump_reverse_0/capacitors_5_0/capacitor_5_3/buffer_and_gate_0/in1 0 2.57f
C413 CP2_5_stage_1/charge_pump_reverse_0/capacitors_5_0/capacitor_5_2/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C414 CP2_5_stage_1/charge_pump_reverse_0/capacitors_5_0/capacitor_5_2/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C415 CP2_5_stage_1/charge_pump_reverse_0/capacitors_5_0/capacitor_5_2/buffer_and_gate_0/in1 0 2.57f
C416 CP2_5_stage_1/charge_pump_reverse_0/capacitors_5_0/capacitor_5_1/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C417 CP2_5_stage_1/charge_pump_reverse_0/capacitors_5_0/capacitor_5_1/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C418 CP2_5_stage_1/charge_pump_reverse_0/capacitors_5_0/capacitor_5_1/buffer_and_gate_0/in1 0 2.57f
C419 CP2_5_stage_1/charge_pump_reverse_0/capacitors_5_0/capacitor_5_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C420 CP2_5_stage_1/charge_pump_reverse_0/capacitors_5_0/capacitor_5_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C421 CP2_5_stage_1/charge_pump_reverse_0/capacitors_5_0/capacitor_5_0/buffer_and_gate_0/in1 0 2.57f
C422 CP2_5_stage_1/charge_pump_reverse_0/nmos_dnw3_0/out1 0 15.1f
C423 CP2_5_stage_1/charge_pump_reverse_0/capacitors_5_0/capacitor_5_7/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C424 CP2_5_stage_1/charge_pump_reverse_0/clock_0/clkb 0 86.4f
C425 CP2_5_stage_1/charge_pump_reverse_0/capacitors_5_0/capacitor_5_7/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C426 CP2_5_stage_1/charge_pump_reverse_0/capacitors_5_0/capacitor_5_7/buffer_and_gate_0/in1 0 2.57f
C427 CP2_5_stage_1/charge_pump_reverse_0/capacitors_5_0/capacitor_5_6/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C428 CP2_5_stage_1/charge_pump_reverse_0/capacitors_5_0/capacitor_5_6/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C429 CP2_5_stage_1/charge_pump_reverse_0/capacitors_5_0/capacitor_5_6/buffer_and_gate_0/in1 0 2.57f
C430 CP2_5_stage_1/charge_pump_reverse_0/capacitors_5_0/capacitor_5_5/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C431 CP2_5_stage_1/charge_pump_reverse_0/capacitors_5_0/capacitor_5_5/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C432 CP2_5_stage_1/charge_pump_reverse_0/capacitors_5_0/capacitor_5_5/buffer_and_gate_0/in1 0 2.57f
C433 CP2_5_stage_1/charge_pump_reverse_0/capacitors_5_1/capacitor_5_4/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C434 CP2_5_stage_1/charge_pump_reverse_0/capacitors_5_1/capacitor_5_4/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C435 CP2_5_stage_1/charge_pump_reverse_0/capacitors_5_1/capacitor_5_4/buffer_and_gate_0/in1 0 2.57f
C436 CP2_5_stage_1/charge_pump_reverse_0/capacitors_5_1/capacitor_5_3/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C437 CP2_5_stage_1/charge_pump_reverse_0/capacitors_5_1/capacitor_5_3/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C438 CP2_5_stage_1/charge_pump_reverse_0/capacitors_5_1/capacitor_5_3/buffer_and_gate_0/in1 0 2.57f
C439 CP2_5_stage_1/charge_pump_reverse_0/capacitors_5_1/capacitor_5_2/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C440 CP2_5_stage_1/charge_pump_reverse_0/capacitors_5_1/capacitor_5_2/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C441 CP2_5_stage_1/charge_pump_reverse_0/capacitors_5_1/capacitor_5_2/buffer_and_gate_0/in1 0 2.57f
C442 CP2_5_stage_1/charge_pump_reverse_0/capacitors_5_1/capacitor_5_1/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C443 CP2_5_stage_1/charge_pump_reverse_0/capacitors_5_1/capacitor_5_1/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C444 CP2_5_stage_1/charge_pump_reverse_0/capacitors_5_1/capacitor_5_1/buffer_and_gate_0/in1 0 2.57f
C445 CP2_5_stage_1/charge_pump_reverse_0/capacitors_5_1/capacitor_5_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C446 CP2_5_stage_1/charge_pump_reverse_0/capacitors_5_1/capacitor_5_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C447 CP2_5_stage_1/charge_pump_reverse_0/capacitors_5_1/capacitor_5_0/buffer_and_gate_0/in1 0 2.57f
C448 CP2_5_stage_1/charge_pump_reverse_0/nmos_dnw3_0/out2 0 14.9f
C449 CP2_5_stage_1/charge_pump_reverse_0/capacitors_5_1/capacitor_5_7/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C450 CP2_5_stage_1/charge_pump_reverse_0/clock_0/clk 0 80f
C451 CP2_5_stage_1/charge_pump_reverse_0/capacitors_5_1/capacitor_5_7/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C452 CP2_5_stage_1/charge_pump_reverse_0/capacitors_5_1/capacitor_5_7/buffer_and_gate_0/in1 0 2.57f
C453 CP2_5_stage_1/charge_pump_reverse_0/capacitors_5_1/capacitor_5_6/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C454 CP2_5_stage_1/charge_pump_reverse_0/capacitors_5_1/capacitor_5_6/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C455 CP2_5_stage_1/charge_pump_reverse_0/capacitors_5_1/capacitor_5_6/buffer_and_gate_0/in1 0 2.57f
C456 CP2_5_stage_1/charge_pump_reverse_0/capacitors_5_1/capacitor_5_5/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C457 CP2_5_stage_1/charge_pump_reverse_0/capacitors_5_1/capacitor_5_5/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C458 CP2_5_stage_1/charge_pump_reverse_0/capacitors_5_1/capacitor_5_5/buffer_and_gate_0/in1 0 2.57f
C459 CP2_5_stage_1/charge_pump_reverse_0/nmos_dnw3_0/clk 0 2.43f
C460 CP2_5_stage_1/m1_94493_n2143# 0 13.9f
C461 CP2_5_stage_1/m1_71529_n2069# 0 3.9f
C462 CP2_5_stage_1/charge_pump_1/clock_0/clk_in 0 13.1f
C463 CP2_5_stage_1/charge_pump_reverse_0/clock_0/clk_in 0 7.77f
C464 CP2_5_stage_1/charge_pump_2/nmos_dnw3_0/vs 0 16.4f
C465 CP2_5_stage_1/charge_pump_2/m1_12174_n760# 0 2.03f
C466 CP2_5_stage_1/charge_pump_2/clock_0/a_2432_n962# 0 8.68f **FLOATING
C467 CP2_5_stage_1/charge_pump_2/clock_0/a_2020_n482# 0 2.57f **FLOATING
C468 CP2_5_stage_1/charge_pump_2/clock_0/a_344_102# 0 2.81f
C469 CP2_5_stage_1/charge_pump_2/clock_0/a_2402_572# 0 2.17f
C470 CP2_5_stage_1/charge_pump_2/clock_0/a_344_n986# 0 2.38f
C471 CP2_5_stage_1/charge_pump_2/clock_0/a_3246_118# 0 6.83f
C472 CP2_5_stage_1/charge_pump_2/nmos_dnw3_0/vin 0 4.17f
C473 CP2_5_stage_1/charge_pump_2/nmos_dnw3_0/clkb 0 2.54f
C474 CP2_5_stage_1/charge_pump_2/capacitors_5_0/capacitor_5_4/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C475 CP2_5_stage_1/charge_pump_2/capacitors_5_0/capacitor_5_4/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C476 CP2_5_stage_1/charge_pump_2/capacitors_5_0/capacitor_5_4/buffer_and_gate_0/in1 0 2.57f
C477 CP2_5_stage_1/charge_pump_2/capacitors_5_0/capacitor_5_3/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C478 CP2_5_stage_1/charge_pump_2/capacitors_5_0/capacitor_5_3/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C479 CP2_5_stage_1/charge_pump_2/capacitors_5_0/capacitor_5_3/buffer_and_gate_0/in1 0 2.57f
C480 CP2_5_stage_1/charge_pump_2/capacitors_5_0/capacitor_5_2/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C481 CP2_5_stage_1/charge_pump_2/capacitors_5_0/capacitor_5_2/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C482 CP2_5_stage_1/charge_pump_2/capacitors_5_0/capacitor_5_2/buffer_and_gate_0/in1 0 2.57f
C483 CP2_5_stage_1/charge_pump_2/capacitors_5_0/capacitor_5_1/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C484 CP2_5_stage_1/charge_pump_2/capacitors_5_0/capacitor_5_1/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C485 CP2_5_stage_1/charge_pump_2/capacitors_5_0/capacitor_5_1/buffer_and_gate_0/in1 0 2.57f
C486 CP2_5_stage_1/charge_pump_2/capacitors_5_0/capacitor_5_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C487 CP2_5_stage_1/charge_pump_2/capacitors_5_0/capacitor_5_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C488 CP2_5_stage_1/charge_pump_2/capacitors_5_0/capacitor_5_0/buffer_and_gate_0/in1 0 2.57f
C489 scanchain_0/data_out[0] 0 37.8f
C490 CP2_5_stage_1/charge_pump_2/nmos_dnw3_0/out1 0 15f
C491 CP2_5_stage_1/charge_pump_2/capacitors_5_0/capacitor_5_7/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C492 CP2_5_stage_1/charge_pump_2/clock_0/clk 0 78.7f
C493 CP2_5_stage_1/charge_pump_2/capacitors_5_0/capacitor_5_7/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C494 CP2_5_stage_1/charge_pump_2/capacitors_5_0/capacitor_5_7/buffer_and_gate_0/in1 0 2.57f
C495 CP2_5_stage_1/charge_pump_2/capacitors_5_0/capacitor_5_6/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C496 CP2_5_stage_1/charge_pump_2/capacitors_5_0/capacitor_5_6/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C497 CP2_5_stage_1/charge_pump_2/capacitors_5_0/capacitor_5_6/buffer_and_gate_0/in1 0 2.57f
C498 CP2_5_stage_1/charge_pump_2/capacitors_5_0/capacitor_5_5/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C499 CP2_5_stage_1/charge_pump_2/capacitors_5_0/capacitor_5_5/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C500 CP2_5_stage_1/charge_pump_2/capacitors_5_0/capacitor_5_5/buffer_and_gate_0/in1 0 2.57f
C501 CP2_5_stage_1/charge_pump_2/capacitors_5_1/capacitor_5_4/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C502 CP2_5_stage_1/charge_pump_2/capacitors_5_1/capacitor_5_4/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C503 CP2_5_stage_1/charge_pump_2/capacitors_5_1/capacitor_5_4/buffer_and_gate_0/in1 0 2.57f
C504 CP2_5_stage_1/charge_pump_2/capacitors_5_1/capacitor_5_3/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C505 CP2_5_stage_1/charge_pump_2/capacitors_5_1/capacitor_5_3/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C506 CP2_5_stage_1/charge_pump_2/capacitors_5_1/capacitor_5_3/buffer_and_gate_0/in1 0 2.57f
C507 CP2_5_stage_1/charge_pump_2/capacitors_5_1/capacitor_5_2/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C508 CP2_5_stage_1/charge_pump_2/capacitors_5_1/capacitor_5_2/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C509 CP2_5_stage_1/charge_pump_2/capacitors_5_1/capacitor_5_2/buffer_and_gate_0/in1 0 2.57f
C510 CP2_5_stage_1/charge_pump_2/capacitors_5_1/capacitor_5_1/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C511 CP2_5_stage_1/charge_pump_2/capacitors_5_1/capacitor_5_1/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C512 CP2_5_stage_1/charge_pump_2/capacitors_5_1/capacitor_5_1/buffer_and_gate_0/in1 0 2.57f
C513 CP2_5_stage_1/charge_pump_2/capacitors_5_1/capacitor_5_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C514 CP2_5_stage_1/charge_pump_2/capacitors_5_1/capacitor_5_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C515 CP2_5_stage_1/charge_pump_2/capacitors_5_1/capacitor_5_0/buffer_and_gate_0/in1 0 2.57f
C516 CP2_5_stage_1/charge_pump_2/nmos_dnw3_0/out2 0 13.6f
C517 CP2_5_stage_1/charge_pump_2/capacitors_5_1/capacitor_5_7/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C518 CP2_5_stage_1/charge_pump_2/clock_0/clkb 0 80.5f
C519 CP2_5_stage_1/charge_pump_2/capacitors_5_1/capacitor_5_7/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C520 CP2_5_stage_1/charge_pump_2/capacitors_5_1/capacitor_5_7/buffer_and_gate_0/in1 0 2.57f
C521 CP2_5_stage_1/charge_pump_2/capacitors_5_1/capacitor_5_6/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C522 CP2_5_stage_1/charge_pump_2/capacitors_5_1/capacitor_5_6/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C523 CP2_5_stage_1/charge_pump_2/capacitors_5_1/capacitor_5_6/buffer_and_gate_0/in1 0 2.57f
C524 CP2_5_stage_1/charge_pump_2/capacitors_5_1/capacitor_5_5/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C525 CP2_5_stage_1/charge_pump_2/capacitors_5_1/capacitor_5_5/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C526 CP2_5_stage_1/charge_pump_2/capacitors_5_1/capacitor_5_5/buffer_and_gate_0/in1 0 2.57f
C527 CP2_5_stage_1/charge_pump_2/nmos_dnw3_0/clk 0 2.76f
C528 CP2_5_stage_1/charge_pump_1/nmos_dnw3_0/vs 0 16.4f
C529 CP2_5_stage_1/charge_pump_reverse_1/nmos_dnw3_0/vin 0 3.91f
C530 CP2_5_stage_1/charge_pump_1/clock_0/a_2432_n962# 0 8.68f **FLOATING
C531 CP2_5_stage_1/charge_pump_1/clock_0/a_2020_n482# 0 2.57f **FLOATING
C532 CP2_5_stage_1/charge_pump_1/clock_0/a_344_102# 0 2.81f
C533 CP2_5_stage_1/charge_pump_1/clock_0/a_2402_572# 0 2.17f
C534 CP2_5_stage_1/charge_pump_1/clock_0/a_344_n986# 0 2.38f
C535 CP2_5_stage_1/charge_pump_1/clock_0/a_3246_118# 0 6.83f
C536 CP2_5_stage_1/charge_pump_1/nmos_dnw3_0/vin 0 4.27f
C537 CP2_5_stage_1/charge_pump_1/nmos_dnw3_0/clkb 0 2.54f
C538 CP2_5_stage_1/charge_pump_1/capacitors_5_0/capacitor_5_4/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C539 CP2_5_stage_1/charge_pump_1/capacitors_5_0/capacitor_5_4/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C540 CP2_5_stage_1/charge_pump_1/capacitors_5_0/capacitor_5_4/buffer_and_gate_0/in1 0 2.57f
C541 scanchain_0/data_out[4] 0 24.3f
C542 CP2_5_stage_1/charge_pump_1/capacitors_5_0/capacitor_5_3/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C543 CP2_5_stage_1/charge_pump_1/capacitors_5_0/capacitor_5_3/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C544 CP2_5_stage_1/charge_pump_1/capacitors_5_0/capacitor_5_3/buffer_and_gate_0/in1 0 2.57f
C545 scanchain_0/data_out[3] 0 23.9f
C546 CP2_5_stage_1/charge_pump_1/capacitors_5_0/capacitor_5_2/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C547 CP2_5_stage_1/charge_pump_1/capacitors_5_0/capacitor_5_2/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C548 CP2_5_stage_1/charge_pump_1/capacitors_5_0/capacitor_5_2/buffer_and_gate_0/in1 0 2.57f
C549 CP2_5_stage_1/charge_pump_1/capacitors_5_0/capacitor_5_1/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C550 CP2_5_stage_1/charge_pump_1/capacitors_5_0/capacitor_5_1/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C551 CP2_5_stage_1/charge_pump_1/capacitors_5_0/capacitor_5_1/buffer_and_gate_0/in1 0 2.57f
C552 CP2_5_stage_1/charge_pump_1/capacitors_5_0/capacitor_5_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C553 CP2_5_stage_1/charge_pump_1/capacitors_5_0/capacitor_5_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C554 CP2_5_stage_1/charge_pump_1/capacitors_5_0/capacitor_5_0/buffer_and_gate_0/in1 0 2.57f
C555 CP2_5_stage_1/charge_pump_1/nmos_dnw3_0/out1 0 15f
C556 CP2_5_stage_1/charge_pump_1/capacitors_5_0/capacitor_5_7/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C557 CP2_5_stage_1/charge_pump_1/clock_0/clk 0 78.7f
C558 CP2_5_stage_1/charge_pump_1/capacitors_5_0/capacitor_5_7/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C559 CP2_5_stage_1/charge_pump_1/capacitors_5_0/capacitor_5_7/buffer_and_gate_0/in1 0 2.57f
C560 scanchain_0/data_out[7] 0 44.5f
C561 CP2_5_stage_1/charge_pump_1/capacitors_5_0/capacitor_5_6/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C562 CP2_5_stage_1/charge_pump_1/capacitors_5_0/capacitor_5_6/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C563 CP2_5_stage_1/charge_pump_1/capacitors_5_0/capacitor_5_6/buffer_and_gate_0/in1 0 2.57f
C564 CP2_5_stage_1/charge_pump_1/capacitors_5_0/capacitor_5_5/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C565 CP2_5_stage_1/charge_pump_1/capacitors_5_0/capacitor_5_5/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C566 CP2_5_stage_1/charge_pump_1/capacitors_5_0/capacitor_5_5/buffer_and_gate_0/in1 0 2.57f
C567 CP2_5_stage_1/charge_pump_1/capacitors_5_1/capacitor_5_4/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C568 CP2_5_stage_1/charge_pump_1/capacitors_5_1/capacitor_5_4/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C569 CP2_5_stage_1/charge_pump_1/capacitors_5_1/capacitor_5_4/buffer_and_gate_0/in1 0 2.57f
C570 CP2_5_stage_1/charge_pump_1/capacitors_5_1/capacitor_5_3/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C571 CP2_5_stage_1/charge_pump_1/capacitors_5_1/capacitor_5_3/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C572 CP2_5_stage_1/charge_pump_1/capacitors_5_1/capacitor_5_3/buffer_and_gate_0/in1 0 2.57f
C573 CP2_5_stage_1/charge_pump_1/capacitors_5_1/capacitor_5_2/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C574 CP2_5_stage_1/charge_pump_1/capacitors_5_1/capacitor_5_2/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C575 CP2_5_stage_1/charge_pump_1/capacitors_5_1/capacitor_5_2/buffer_and_gate_0/in1 0 2.57f
C576 CP2_5_stage_1/charge_pump_1/capacitors_5_1/capacitor_5_1/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C577 CP2_5_stage_1/charge_pump_1/capacitors_5_1/capacitor_5_1/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C578 CP2_5_stage_1/charge_pump_1/capacitors_5_1/capacitor_5_1/buffer_and_gate_0/in1 0 2.57f
C579 CP2_5_stage_1/charge_pump_1/capacitors_5_1/capacitor_5_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C580 CP2_5_stage_1/charge_pump_1/capacitors_5_1/capacitor_5_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C581 CP2_5_stage_1/charge_pump_1/capacitors_5_1/capacitor_5_0/buffer_and_gate_0/in1 0 2.57f
C582 CP2_5_stage_1/charge_pump_1/nmos_dnw3_0/out2 0 13.6f
C583 CP2_5_stage_1/charge_pump_1/capacitors_5_1/capacitor_5_7/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C584 CP2_5_stage_1/charge_pump_1/clock_0/clkb 0 80.5f
C585 CP2_5_stage_1/charge_pump_1/capacitors_5_1/capacitor_5_7/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C586 CP2_5_stage_1/charge_pump_1/capacitors_5_1/capacitor_5_7/buffer_and_gate_0/in1 0 2.57f
C587 CP2_5_stage_1/charge_pump_1/capacitors_5_1/capacitor_5_6/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C588 CP2_5_stage_1/charge_pump_1/capacitors_5_1/capacitor_5_6/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C589 CP2_5_stage_1/charge_pump_1/capacitors_5_1/capacitor_5_6/buffer_and_gate_0/in1 0 2.57f
C590 CP2_5_stage_1/charge_pump_1/capacitors_5_1/capacitor_5_5/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C591 CP2_5_stage_1/charge_pump_1/capacitors_5_1/capacitor_5_5/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C592 CP2_5_stage_1/charge_pump_1/capacitors_5_1/capacitor_5_5/buffer_and_gate_0/in1 0 2.57f
C593 CP2_5_stage_1/charge_pump_1/nmos_dnw3_0/clk 0 2.76f
C594 CP2_5_stage_1/charge_pump_0/nmos_dnw3_0/vs 0 16.4f
C595 CP2_5_stage_1/charge_pump_reverse_0/nmos_dnw3_0/vin 0 2.33f
C596 CP2_5_stage_1/charge_pump_0/clock_0/a_2432_n962# 0 8.68f **FLOATING
C597 CP2_5_stage_1/charge_pump_0/clock_0/a_2020_n482# 0 2.57f **FLOATING
C598 CP2_5_stage_1/charge_pump_0/clock_0/a_344_102# 0 2.81f
C599 CP2_5_stage_1/charge_pump_0/clock_0/a_2402_572# 0 2.17f
C600 CP2_5_stage_1/charge_pump_0/clock_0/a_344_n986# 0 2.38f
C601 CP1_5_stage_0/charge_pump1_0/clk_in 0 91.3f
C602 CP2_5_stage_1/charge_pump_0/clock_0/a_3246_118# 0 6.83f
C603 CP2_5_stage_1/charge_pump_0/nmos_dnw3_0/vin 0 2.94f
C604 CP2_5_stage_1/charge_pump_0/nmos_dnw3_0/clkb 0 2.54f
C605 CP2_5_stage_1/charge_pump_0/capacitors_5_0/capacitor_5_4/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C606 CP2_5_stage_1/charge_pump_0/capacitors_5_0/capacitor_5_4/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C607 CP2_5_stage_1/charge_pump_0/capacitors_5_0/capacitor_5_4/buffer_and_gate_0/in1 0 2.57f
C608 CP2_5_stage_1/charge_pump_0/capacitors_5_0/capacitor_5_3/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C609 CP2_5_stage_1/charge_pump_0/capacitors_5_0/capacitor_5_3/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C610 CP2_5_stage_1/charge_pump_0/capacitors_5_0/capacitor_5_3/buffer_and_gate_0/in1 0 2.57f
C611 CP2_5_stage_1/charge_pump_0/capacitors_5_0/capacitor_5_2/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C612 CP2_5_stage_1/charge_pump_0/capacitors_5_0/capacitor_5_2/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C613 CP2_5_stage_1/charge_pump_0/capacitors_5_0/capacitor_5_2/buffer_and_gate_0/in1 0 2.57f
C614 CP2_5_stage_1/charge_pump_0/capacitors_5_0/capacitor_5_1/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C615 CP2_5_stage_1/charge_pump_0/capacitors_5_0/capacitor_5_1/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C616 CP2_5_stage_1/charge_pump_0/capacitors_5_0/capacitor_5_1/buffer_and_gate_0/in1 0 2.57f
C617 CP2_5_stage_1/charge_pump_0/capacitors_5_0/capacitor_5_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C618 CP2_5_stage_1/charge_pump_0/capacitors_5_0/capacitor_5_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C619 CP2_5_stage_1/charge_pump_0/capacitors_5_0/capacitor_5_0/buffer_and_gate_0/in1 0 2.57f
C620 CP2_5_stage_1/charge_pump_0/nmos_dnw3_0/out1 0 15f
C621 CP2_5_stage_1/charge_pump_0/capacitors_5_0/capacitor_5_7/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C622 CP2_5_stage_1/charge_pump_0/clock_0/clk 0 78.7f
C623 CP2_5_stage_1/charge_pump_0/capacitors_5_0/capacitor_5_7/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C624 VSUBS 0 1.82p
C625 CP2_5_stage_1/charge_pump_0/capacitors_5_0/capacitor_5_7/buffer_and_gate_0/in1 0 2.57f
C626 CP2_5_stage_1/charge_pump_0/capacitors_5_0/capacitor_5_6/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C627 CP2_5_stage_1/charge_pump_0/capacitors_5_0/capacitor_5_6/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C628 CP2_5_stage_1/charge_pump_0/capacitors_5_0/capacitor_5_6/buffer_and_gate_0/in1 0 2.57f
C629 scanchain_0/data_out[6] 0 41.6f
C630 CP2_5_stage_1/charge_pump_0/capacitors_5_0/capacitor_5_5/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C631 CP2_5_stage_1/charge_pump_0/capacitors_5_0/capacitor_5_5/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C632 CP2_5_stage_1/charge_pump_0/capacitors_5_0/capacitor_5_5/buffer_and_gate_0/in1 0 2.57f
C633 scanchain_0/data_out[5] 0 32.3f
C634 CP2_5_stage_1/charge_pump_0/capacitors_5_1/capacitor_5_4/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C635 CP2_5_stage_1/charge_pump_0/capacitors_5_1/capacitor_5_4/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C636 CP2_5_stage_1/charge_pump_0/capacitors_5_1/capacitor_5_4/buffer_and_gate_0/in1 0 2.57f
C637 CP2_5_stage_1/charge_pump_0/capacitors_5_1/capacitor_5_3/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C638 CP2_5_stage_1/charge_pump_0/capacitors_5_1/capacitor_5_3/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C639 CP2_5_stage_1/charge_pump_0/capacitors_5_1/capacitor_5_3/buffer_and_gate_0/in1 0 2.57f
C640 CP2_5_stage_1/charge_pump_0/capacitors_5_1/capacitor_5_2/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C641 CP2_5_stage_1/charge_pump_0/capacitors_5_1/capacitor_5_2/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C642 CP2_5_stage_1/charge_pump_0/capacitors_5_1/capacitor_5_2/buffer_and_gate_0/in1 0 2.57f
C643 CP2_5_stage_1/charge_pump_0/capacitors_5_1/capacitor_5_1/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C644 CP2_5_stage_1/charge_pump_0/capacitors_5_1/capacitor_5_1/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C645 CP2_5_stage_1/charge_pump_0/capacitors_5_1/capacitor_5_1/buffer_and_gate_0/in1 0 2.57f
C646 CP2_5_stage_1/charge_pump_0/capacitors_5_1/capacitor_5_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C647 CP2_5_stage_1/charge_pump_0/capacitors_5_1/capacitor_5_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C648 CP2_5_stage_1/charge_pump_0/capacitors_5_1/capacitor_5_0/buffer_and_gate_0/in1 0 2.57f
C649 CP2_5_stage_1/charge_pump_0/nmos_dnw3_0/out2 0 13.6f
C650 CP2_5_stage_1/charge_pump_0/capacitors_5_1/capacitor_5_7/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C651 CP2_5_stage_1/charge_pump_0/clock_0/clkb 0 80.5f
C652 CP2_5_stage_1/charge_pump_0/capacitors_5_1/capacitor_5_7/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C653 CP1_5_stage_0/charge_pump1_2/vdd 0 7.22p
C654 CP2_5_stage_1/charge_pump_0/capacitors_5_1/capacitor_5_7/buffer_and_gate_0/in1 0 2.57f
C655 CP2_5_stage_1/charge_pump_0/capacitors_5_1/capacitor_5_6/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C656 CP2_5_stage_1/charge_pump_0/capacitors_5_1/capacitor_5_6/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C657 CP2_5_stage_1/charge_pump_0/capacitors_5_1/capacitor_5_6/buffer_and_gate_0/in1 0 2.57f
C658 CP2_5_stage_1/charge_pump_0/capacitors_5_1/capacitor_5_5/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C659 CP2_5_stage_1/charge_pump_0/capacitors_5_1/capacitor_5_5/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C660 CP2_5_stage_1/charge_pump_0/capacitors_5_1/capacitor_5_5/buffer_and_gate_0/in1 0 2.57f
C661 CP2_5_stage_1/charge_pump_0/nmos_dnw3_0/clk 0 2.76f
C662 CP2_5_stage_0/charge_pump_reverse_1/nmos_dnw3_0/vs 0 16.4f
C663 CP2_5_stage_0/charge_pump_reverse_1/sky130_fd_pr__pfet_01v8_4RPJ49_1/w_n3905_n142# 0 6.63f
C664 CP2_5_stage_0/charge_pump_reverse_1/sky130_fd_pr__pfet_01v8_4RPJ49_0/w_n3905_n142# 0 6.63f
C665 CP2_5_stage_0/charge_pump_reverse_1/clock_0/a_2432_n962# 0 8.68f **FLOATING
C666 CP2_5_stage_0/charge_pump_reverse_1/clock_0/a_2020_n482# 0 2.57f **FLOATING
C667 CP2_5_stage_0/charge_pump_reverse_1/clock_0/a_344_102# 0 2.81f
C668 CP2_5_stage_0/charge_pump_reverse_1/clock_0/a_2402_572# 0 2.17f
C669 CP2_5_stage_0/charge_pump_reverse_1/clock_0/a_344_n986# 0 2.38f
C670 CP2_5_stage_0/charge_pump_reverse_1/clock_0/a_3246_118# 0 6.83f
C671 CP2_5_stage_0/charge_pump_reverse_1/nmos_dnw3_0/clkb 0 2.23f
C672 CP2_5_stage_0/charge_pump_reverse_1/capacitors_5_0/capacitor_5_4/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C673 CP2_5_stage_0/charge_pump_reverse_1/capacitors_5_0/capacitor_5_4/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C674 CP2_5_stage_0/charge_pump_reverse_1/capacitors_5_0/capacitor_5_4/buffer_and_gate_0/in1 0 2.57f
C675 CP2_5_stage_0/charge_pump_reverse_1/capacitors_5_0/capacitor_5_3/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C676 CP2_5_stage_0/charge_pump_reverse_1/capacitors_5_0/capacitor_5_3/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C677 CP2_5_stage_0/charge_pump_reverse_1/capacitors_5_0/capacitor_5_3/buffer_and_gate_0/in1 0 2.57f
C678 CP2_5_stage_0/charge_pump_reverse_1/capacitors_5_0/capacitor_5_2/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C679 CP2_5_stage_0/charge_pump_reverse_1/capacitors_5_0/capacitor_5_2/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C680 CP2_5_stage_0/charge_pump_reverse_1/capacitors_5_0/capacitor_5_2/buffer_and_gate_0/in1 0 2.57f
C681 CP2_5_stage_0/charge_pump_reverse_1/capacitors_5_0/capacitor_5_1/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C682 CP2_5_stage_0/charge_pump_reverse_1/capacitors_5_0/capacitor_5_1/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C683 CP2_5_stage_0/charge_pump_reverse_1/capacitors_5_0/capacitor_5_1/buffer_and_gate_0/in1 0 2.57f
C684 CP2_5_stage_0/charge_pump_reverse_1/capacitors_5_0/capacitor_5_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C685 CP2_5_stage_0/charge_pump_reverse_1/capacitors_5_0/capacitor_5_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C686 CP2_5_stage_0/charge_pump_reverse_1/capacitors_5_0/capacitor_5_0/buffer_and_gate_0/in1 0 2.57f
C687 CP2_5_stage_0/charge_pump_reverse_1/nmos_dnw3_0/out1 0 15.1f
C688 CP2_5_stage_0/charge_pump_reverse_1/capacitors_5_0/capacitor_5_7/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C689 CP2_5_stage_0/charge_pump_reverse_1/clock_0/clkb 0 86.4f
C690 CP2_5_stage_0/charge_pump_reverse_1/capacitors_5_0/capacitor_5_7/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C691 CP2_5_stage_0/charge_pump_reverse_1/capacitors_5_0/capacitor_5_7/buffer_and_gate_0/in1 0 2.57f
C692 CP2_5_stage_0/charge_pump_reverse_1/capacitors_5_0/capacitor_5_6/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C693 CP2_5_stage_0/charge_pump_reverse_1/capacitors_5_0/capacitor_5_6/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C694 CP2_5_stage_0/charge_pump_reverse_1/capacitors_5_0/capacitor_5_6/buffer_and_gate_0/in1 0 2.57f
C695 CP2_5_stage_0/charge_pump_reverse_1/capacitors_5_0/capacitor_5_5/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C696 CP2_5_stage_0/charge_pump_reverse_1/capacitors_5_0/capacitor_5_5/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C697 CP2_5_stage_0/charge_pump_reverse_1/capacitors_5_0/capacitor_5_5/buffer_and_gate_0/in1 0 2.57f
C698 CP2_5_stage_0/charge_pump_reverse_1/capacitors_5_1/capacitor_5_4/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C699 CP2_5_stage_0/charge_pump_reverse_1/capacitors_5_1/capacitor_5_4/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C700 CP2_5_stage_0/charge_pump_reverse_1/capacitors_5_1/capacitor_5_4/buffer_and_gate_0/in1 0 2.57f
C701 CP2_5_stage_0/charge_pump_reverse_1/capacitors_5_1/capacitor_5_3/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C702 CP2_5_stage_0/charge_pump_reverse_1/capacitors_5_1/capacitor_5_3/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C703 CP2_5_stage_0/charge_pump_reverse_1/capacitors_5_1/capacitor_5_3/buffer_and_gate_0/in1 0 2.57f
C704 CP2_5_stage_0/charge_pump_reverse_1/capacitors_5_1/capacitor_5_2/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C705 CP2_5_stage_0/charge_pump_reverse_1/capacitors_5_1/capacitor_5_2/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C706 CP2_5_stage_0/charge_pump_reverse_1/capacitors_5_1/capacitor_5_2/buffer_and_gate_0/in1 0 2.57f
C707 CP2_5_stage_0/charge_pump_reverse_1/capacitors_5_1/capacitor_5_1/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C708 CP2_5_stage_0/charge_pump_reverse_1/capacitors_5_1/capacitor_5_1/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C709 CP2_5_stage_0/charge_pump_reverse_1/capacitors_5_1/capacitor_5_1/buffer_and_gate_0/in1 0 2.57f
C710 CP2_5_stage_0/charge_pump_reverse_1/capacitors_5_1/capacitor_5_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C711 CP2_5_stage_0/charge_pump_reverse_1/capacitors_5_1/capacitor_5_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C712 CP2_5_stage_0/charge_pump_reverse_1/capacitors_5_1/capacitor_5_0/buffer_and_gate_0/in1 0 2.57f
C713 CP2_5_stage_0/charge_pump_reverse_1/capacitors_5_1/capacitor_5_7/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C714 CP2_5_stage_0/charge_pump_reverse_1/capacitors_5_1/capacitor_5_7/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C715 CP2_5_stage_0/charge_pump_reverse_1/capacitors_5_1/capacitor_5_7/buffer_and_gate_0/in1 0 2.57f
C716 CP2_5_stage_0/charge_pump_reverse_1/capacitors_5_1/capacitor_5_6/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C717 CP2_5_stage_0/charge_pump_reverse_1/capacitors_5_1/capacitor_5_6/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C718 CP2_5_stage_0/charge_pump_reverse_1/capacitors_5_1/capacitor_5_6/buffer_and_gate_0/in1 0 2.57f
C719 CP2_5_stage_0/charge_pump_reverse_1/capacitors_5_1/capacitor_5_5/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C720 CP2_5_stage_0/charge_pump_reverse_1/capacitors_5_1/capacitor_5_5/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C721 CP2_5_stage_0/charge_pump_reverse_1/capacitors_5_1/capacitor_5_5/buffer_and_gate_0/in1 0 2.57f
C722 CP2_5_stage_0/charge_pump_reverse_1/nmos_dnw3_0/clk 0 2.43f
C723 CP2_5_stage_0/charge_pump_reverse_0/nmos_dnw3_0/vs 0 16.4f
C724 CP2_5_stage_0/charge_pump_reverse_0/sky130_fd_pr__pfet_01v8_4RPJ49_1/w_n3905_n142# 0 6.63f
C725 CP2_5_stage_0/charge_pump_reverse_0/sky130_fd_pr__pfet_01v8_4RPJ49_0/w_n3905_n142# 0 6.63f
C726 CP2_5_stage_0/charge_pump_reverse_0/clock_0/a_2432_n962# 0 8.68f **FLOATING
C727 CP2_5_stage_0/charge_pump_reverse_0/clock_0/a_2020_n482# 0 2.57f **FLOATING
C728 CP2_5_stage_0/charge_pump_reverse_0/clock_0/a_344_102# 0 2.81f
C729 CP2_5_stage_0/charge_pump_reverse_0/clock_0/a_2402_572# 0 2.17f
C730 CP2_5_stage_0/charge_pump_reverse_0/clock_0/a_344_n986# 0 2.38f
C731 CP2_5_stage_0/charge_pump_reverse_0/clock_0/a_3246_118# 0 6.83f
C732 CP2_5_stage_0/charge_pump_reverse_0/nmos_dnw3_0/clkb 0 2.23f
C733 CP2_5_stage_0/charge_pump_reverse_0/capacitors_5_0/capacitor_5_4/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C734 CP2_5_stage_0/charge_pump_reverse_0/capacitors_5_0/capacitor_5_4/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C735 CP2_5_stage_0/charge_pump_reverse_0/capacitors_5_0/capacitor_5_4/buffer_and_gate_0/in1 0 2.57f
C736 CP2_5_stage_0/charge_pump_reverse_0/capacitors_5_0/capacitor_5_3/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C737 CP2_5_stage_0/charge_pump_reverse_0/capacitors_5_0/capacitor_5_3/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C738 CP2_5_stage_0/charge_pump_reverse_0/capacitors_5_0/capacitor_5_3/buffer_and_gate_0/in1 0 2.57f
C739 CP2_5_stage_0/charge_pump_reverse_0/capacitors_5_0/capacitor_5_2/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C740 CP2_5_stage_0/charge_pump_reverse_0/capacitors_5_0/capacitor_5_2/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C741 CP2_5_stage_0/charge_pump_reverse_0/capacitors_5_0/capacitor_5_2/buffer_and_gate_0/in1 0 2.57f
C742 CP2_5_stage_0/charge_pump_reverse_0/capacitors_5_0/capacitor_5_1/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C743 CP2_5_stage_0/charge_pump_reverse_0/capacitors_5_0/capacitor_5_1/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C744 CP2_5_stage_0/charge_pump_reverse_0/capacitors_5_0/capacitor_5_1/buffer_and_gate_0/in1 0 2.57f
C745 CP2_5_stage_0/charge_pump_reverse_0/capacitors_5_0/capacitor_5_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C746 CP2_5_stage_0/charge_pump_reverse_0/capacitors_5_0/capacitor_5_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C747 CP2_5_stage_0/charge_pump_reverse_0/capacitors_5_0/capacitor_5_0/buffer_and_gate_0/in1 0 2.57f
C748 CP2_5_stage_0/charge_pump_reverse_0/nmos_dnw3_0/out1 0 15.1f
C749 CP2_5_stage_0/charge_pump_reverse_0/capacitors_5_0/capacitor_5_7/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C750 CP2_5_stage_0/charge_pump_reverse_0/clock_0/clkb 0 86.4f
C751 CP2_5_stage_0/charge_pump_reverse_0/capacitors_5_0/capacitor_5_7/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C752 CP2_5_stage_0/charge_pump_reverse_0/capacitors_5_0/capacitor_5_7/buffer_and_gate_0/in1 0 2.57f
C753 CP2_5_stage_0/charge_pump_reverse_0/capacitors_5_0/capacitor_5_6/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C754 CP2_5_stage_0/charge_pump_reverse_0/capacitors_5_0/capacitor_5_6/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C755 CP2_5_stage_0/charge_pump_reverse_0/capacitors_5_0/capacitor_5_6/buffer_and_gate_0/in1 0 2.57f
C756 CP2_5_stage_0/charge_pump_reverse_0/capacitors_5_0/capacitor_5_5/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C757 CP2_5_stage_0/charge_pump_reverse_0/capacitors_5_0/capacitor_5_5/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C758 CP2_5_stage_0/charge_pump_reverse_0/capacitors_5_0/capacitor_5_5/buffer_and_gate_0/in1 0 2.57f
C759 CP2_5_stage_0/charge_pump_reverse_0/capacitors_5_1/capacitor_5_4/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C760 CP2_5_stage_0/charge_pump_reverse_0/capacitors_5_1/capacitor_5_4/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C761 CP2_5_stage_0/charge_pump_reverse_0/capacitors_5_1/capacitor_5_4/buffer_and_gate_0/in1 0 2.57f
C762 CP2_5_stage_0/charge_pump_reverse_0/capacitors_5_1/capacitor_5_3/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C763 CP2_5_stage_0/charge_pump_reverse_0/capacitors_5_1/capacitor_5_3/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C764 CP2_5_stage_0/charge_pump_reverse_0/capacitors_5_1/capacitor_5_3/buffer_and_gate_0/in1 0 2.57f
C765 CP2_5_stage_0/charge_pump_reverse_0/capacitors_5_1/capacitor_5_2/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C766 CP2_5_stage_0/charge_pump_reverse_0/capacitors_5_1/capacitor_5_2/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C767 CP2_5_stage_0/charge_pump_reverse_0/capacitors_5_1/capacitor_5_2/buffer_and_gate_0/in1 0 2.57f
C768 CP2_5_stage_0/charge_pump_reverse_0/capacitors_5_1/capacitor_5_1/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C769 CP2_5_stage_0/charge_pump_reverse_0/capacitors_5_1/capacitor_5_1/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C770 CP2_5_stage_0/charge_pump_reverse_0/capacitors_5_1/capacitor_5_1/buffer_and_gate_0/in1 0 2.57f
C771 CP2_5_stage_0/charge_pump_reverse_0/capacitors_5_1/capacitor_5_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C772 CP2_5_stage_0/charge_pump_reverse_0/capacitors_5_1/capacitor_5_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C773 CP2_5_stage_0/charge_pump_reverse_0/capacitors_5_1/capacitor_5_0/buffer_and_gate_0/in1 0 2.57f
C774 CP2_5_stage_0/charge_pump_reverse_0/nmos_dnw3_0/out2 0 14.9f
C775 CP2_5_stage_0/charge_pump_reverse_0/capacitors_5_1/capacitor_5_7/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C776 CP2_5_stage_0/charge_pump_reverse_0/clock_0/clk 0 80f
C777 CP2_5_stage_0/charge_pump_reverse_0/capacitors_5_1/capacitor_5_7/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C778 CP2_5_stage_0/charge_pump_reverse_0/capacitors_5_1/capacitor_5_7/buffer_and_gate_0/in1 0 2.57f
C779 CP2_5_stage_0/charge_pump_reverse_0/capacitors_5_1/capacitor_5_6/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C780 CP2_5_stage_0/charge_pump_reverse_0/capacitors_5_1/capacitor_5_6/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C781 CP2_5_stage_0/charge_pump_reverse_0/capacitors_5_1/capacitor_5_6/buffer_and_gate_0/in1 0 2.57f
C782 CP2_5_stage_0/charge_pump_reverse_0/capacitors_5_1/capacitor_5_5/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C783 CP2_5_stage_0/charge_pump_reverse_0/capacitors_5_1/capacitor_5_5/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C784 CP2_5_stage_0/charge_pump_reverse_0/capacitors_5_1/capacitor_5_5/buffer_and_gate_0/in1 0 2.57f
C785 CP2_5_stage_0/charge_pump_reverse_0/nmos_dnw3_0/clk 0 2.43f
C786 CP2_5_stage_0/charge_pump_reverse_1/clock_0/clk_in 0 5.88f
C787 CP2_5_stage_0/charge_pump_1/clock_0/clk_in 0 13.1f
C788 CP2_5_stage_0/charge_pump_reverse_0/clock_0/clk_in 0 7.77f
C789 CP2_5_stage_0/charge_pump_2/nmos_dnw3_0/vs 0 16.4f
C790 CP2_5_stage_0/charge_pump_2/clock_0/a_2432_n962# 0 8.68f **FLOATING
C791 CP2_5_stage_0/charge_pump_2/clock_0/a_2020_n482# 0 2.57f **FLOATING
C792 CP2_5_stage_0/charge_pump_2/clock_0/a_344_102# 0 2.81f
C793 CP2_5_stage_0/charge_pump_2/clock_0/a_2402_572# 0 2.17f
C794 CP2_5_stage_0/charge_pump_2/clock_0/a_344_n986# 0 2.38f
C795 CP2_5_stage_0/charge_pump_2/clock_0/a_3246_118# 0 6.83f
C796 CP2_5_stage_0/charge_pump_2/nmos_dnw3_0/vin 0 4.17f
C797 CP2_5_stage_0/charge_pump_2/nmos_dnw3_0/clkb 0 2.54f
C798 CP2_5_stage_0/charge_pump_2/capacitors_5_0/capacitor_5_4/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C799 CP2_5_stage_0/charge_pump_2/capacitors_5_0/capacitor_5_4/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C800 CP2_5_stage_0/charge_pump_2/capacitors_5_0/capacitor_5_4/buffer_and_gate_0/in1 0 2.57f
C801 CP2_5_stage_0/charge_pump_2/capacitors_5_0/capacitor_5_3/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C802 CP2_5_stage_0/charge_pump_2/capacitors_5_0/capacitor_5_3/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C803 CP2_5_stage_0/charge_pump_2/capacitors_5_0/capacitor_5_3/buffer_and_gate_0/in1 0 2.57f
C804 CP2_5_stage_0/charge_pump_2/capacitors_5_0/capacitor_5_2/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C805 CP2_5_stage_0/charge_pump_2/capacitors_5_0/capacitor_5_2/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C806 CP2_5_stage_0/charge_pump_2/capacitors_5_0/capacitor_5_2/buffer_and_gate_0/in1 0 2.57f
C807 CP2_5_stage_0/charge_pump_2/capacitors_5_0/capacitor_5_1/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C808 CP2_5_stage_0/charge_pump_2/capacitors_5_0/capacitor_5_1/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C809 CP2_5_stage_0/charge_pump_2/capacitors_5_0/capacitor_5_1/buffer_and_gate_0/in1 0 2.57f
C810 CP2_5_stage_0/charge_pump_2/capacitors_5_0/capacitor_5_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C811 CP2_5_stage_0/charge_pump_2/capacitors_5_0/capacitor_5_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C812 CP2_5_stage_0/charge_pump_2/capacitors_5_0/capacitor_5_0/buffer_and_gate_0/in1 0 2.57f
C813 CP2_5_stage_0/charge_pump_2/nmos_dnw3_0/out1 0 15f
C814 CP2_5_stage_0/charge_pump_2/capacitors_5_0/capacitor_5_7/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C815 CP2_5_stage_0/charge_pump_2/clock_0/clk 0 78.7f
C816 CP2_5_stage_0/charge_pump_2/capacitors_5_0/capacitor_5_7/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C817 CP2_5_stage_0/charge_pump_2/capacitors_5_0/capacitor_5_7/buffer_and_gate_0/in1 0 2.57f
C818 CP2_5_stage_0/charge_pump_2/capacitors_5_0/capacitor_5_6/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C819 CP2_5_stage_0/charge_pump_2/capacitors_5_0/capacitor_5_6/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C820 CP2_5_stage_0/charge_pump_2/capacitors_5_0/capacitor_5_6/buffer_and_gate_0/in1 0 2.57f
C821 CP2_5_stage_0/charge_pump_2/capacitors_5_0/capacitor_5_5/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C822 CP2_5_stage_0/charge_pump_2/capacitors_5_0/capacitor_5_5/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C823 CP2_5_stage_0/charge_pump_2/capacitors_5_0/capacitor_5_5/buffer_and_gate_0/in1 0 2.57f
C824 CP2_5_stage_0/charge_pump_2/capacitors_5_1/capacitor_5_4/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C825 CP2_5_stage_0/charge_pump_2/capacitors_5_1/capacitor_5_4/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C826 CP2_5_stage_0/charge_pump_2/capacitors_5_1/capacitor_5_4/buffer_and_gate_0/in1 0 2.57f
C827 CP2_5_stage_0/charge_pump_2/capacitors_5_1/capacitor_5_3/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C828 CP2_5_stage_0/charge_pump_2/capacitors_5_1/capacitor_5_3/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C829 CP2_5_stage_0/charge_pump_2/capacitors_5_1/capacitor_5_3/buffer_and_gate_0/in1 0 2.57f
C830 CP2_5_stage_0/charge_pump_2/capacitors_5_1/capacitor_5_2/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C831 CP2_5_stage_0/charge_pump_2/capacitors_5_1/capacitor_5_2/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C832 CP2_5_stage_0/charge_pump_2/capacitors_5_1/capacitor_5_2/buffer_and_gate_0/in1 0 2.57f
C833 CP2_5_stage_0/charge_pump_2/capacitors_5_1/capacitor_5_1/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C834 CP2_5_stage_0/charge_pump_2/capacitors_5_1/capacitor_5_1/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C835 CP2_5_stage_0/charge_pump_2/capacitors_5_1/capacitor_5_1/buffer_and_gate_0/in1 0 2.57f
C836 CP2_5_stage_0/charge_pump_2/capacitors_5_1/capacitor_5_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C837 CP2_5_stage_0/charge_pump_2/capacitors_5_1/capacitor_5_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C838 CP2_5_stage_0/charge_pump_2/capacitors_5_1/capacitor_5_0/buffer_and_gate_0/in1 0 2.57f
C839 CP2_5_stage_0/charge_pump_2/nmos_dnw3_0/out2 0 13.6f
C840 CP2_5_stage_0/charge_pump_2/capacitors_5_1/capacitor_5_7/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C841 CP2_5_stage_0/charge_pump_2/clock_0/clkb 0 80.5f
C842 CP2_5_stage_0/charge_pump_2/capacitors_5_1/capacitor_5_7/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C843 CP2_5_stage_0/charge_pump_2/capacitors_5_1/capacitor_5_7/buffer_and_gate_0/in1 0 2.57f
C844 CP2_5_stage_0/charge_pump_2/capacitors_5_1/capacitor_5_6/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C845 CP2_5_stage_0/charge_pump_2/capacitors_5_1/capacitor_5_6/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C846 CP2_5_stage_0/charge_pump_2/capacitors_5_1/capacitor_5_6/buffer_and_gate_0/in1 0 2.57f
C847 CP2_5_stage_0/charge_pump_2/capacitors_5_1/capacitor_5_5/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C848 CP2_5_stage_0/charge_pump_2/capacitors_5_1/capacitor_5_5/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C849 CP2_5_stage_0/charge_pump_2/capacitors_5_1/capacitor_5_5/buffer_and_gate_0/in1 0 2.57f
C850 CP2_5_stage_0/charge_pump_2/nmos_dnw3_0/clk 0 2.76f
C851 CP2_5_stage_0/charge_pump_1/nmos_dnw3_0/vs 0 16.4f
C852 CP2_5_stage_0/charge_pump_reverse_1/nmos_dnw3_0/vin 0 3.91f
C853 CP2_5_stage_0/charge_pump_1/clock_0/a_2432_n962# 0 8.68f **FLOATING
C854 CP2_5_stage_0/charge_pump_1/clock_0/a_2020_n482# 0 2.57f **FLOATING
C855 CP2_5_stage_0/charge_pump_1/clock_0/a_344_102# 0 2.81f
C856 CP2_5_stage_0/charge_pump_1/clock_0/a_2402_572# 0 2.17f
C857 CP2_5_stage_0/charge_pump_1/clock_0/a_344_n986# 0 2.38f
C858 CP2_5_stage_0/charge_pump_1/clock_0/a_3246_118# 0 6.83f
C859 CP2_5_stage_0/charge_pump_1/nmos_dnw3_0/vin 0 4.27f
C860 CP2_5_stage_0/charge_pump_1/nmos_dnw3_0/clkb 0 2.54f
C861 CP2_5_stage_0/charge_pump_1/capacitors_5_0/capacitor_5_4/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C862 CP2_5_stage_0/charge_pump_1/capacitors_5_0/capacitor_5_4/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C863 CP2_5_stage_0/charge_pump_1/capacitors_5_0/capacitor_5_4/buffer_and_gate_0/in1 0 2.57f
C864 CP2_5_stage_0/charge_pump_1/capacitors_5_0/capacitor_5_3/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C865 CP2_5_stage_0/charge_pump_1/capacitors_5_0/capacitor_5_3/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C866 CP2_5_stage_0/charge_pump_1/capacitors_5_0/capacitor_5_3/buffer_and_gate_0/in1 0 2.57f
C867 CP2_5_stage_0/charge_pump_1/capacitors_5_0/capacitor_5_2/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C868 CP2_5_stage_0/charge_pump_1/capacitors_5_0/capacitor_5_2/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C869 CP2_5_stage_0/charge_pump_1/capacitors_5_0/capacitor_5_2/buffer_and_gate_0/in1 0 2.57f
C870 CP2_5_stage_0/charge_pump_1/capacitors_5_0/capacitor_5_1/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C871 CP2_5_stage_0/charge_pump_1/capacitors_5_0/capacitor_5_1/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C872 CP2_5_stage_0/charge_pump_1/capacitors_5_0/capacitor_5_1/buffer_and_gate_0/in1 0 2.57f
C873 CP2_5_stage_0/charge_pump_1/capacitors_5_0/capacitor_5_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C874 CP2_5_stage_0/charge_pump_1/capacitors_5_0/capacitor_5_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C875 CP2_5_stage_0/charge_pump_1/capacitors_5_0/capacitor_5_0/buffer_and_gate_0/in1 0 2.57f
C876 CP2_5_stage_0/charge_pump_1/nmos_dnw3_0/out1 0 15f
C877 CP2_5_stage_0/charge_pump_1/capacitors_5_0/capacitor_5_7/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C878 CP2_5_stage_0/charge_pump_1/clock_0/clk 0 78.7f
C879 CP2_5_stage_0/charge_pump_1/capacitors_5_0/capacitor_5_7/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C880 CP2_5_stage_0/charge_pump_1/capacitors_5_0/capacitor_5_7/buffer_and_gate_0/in1 0 2.57f
C881 CP2_5_stage_0/charge_pump_1/capacitors_5_0/capacitor_5_6/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C882 CP2_5_stage_0/charge_pump_1/capacitors_5_0/capacitor_5_6/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C883 CP2_5_stage_0/charge_pump_1/capacitors_5_0/capacitor_5_6/buffer_and_gate_0/in1 0 2.57f
C884 CP2_5_stage_0/charge_pump_1/capacitors_5_0/capacitor_5_5/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C885 CP2_5_stage_0/charge_pump_1/capacitors_5_0/capacitor_5_5/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C886 CP2_5_stage_0/charge_pump_1/capacitors_5_0/capacitor_5_5/buffer_and_gate_0/in1 0 2.57f
C887 CP2_5_stage_0/charge_pump_1/capacitors_5_1/capacitor_5_4/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C888 CP2_5_stage_0/charge_pump_1/capacitors_5_1/capacitor_5_4/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C889 CP2_5_stage_0/charge_pump_1/capacitors_5_1/capacitor_5_4/buffer_and_gate_0/in1 0 2.57f
C890 CP2_5_stage_0/charge_pump_1/capacitors_5_1/capacitor_5_3/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C891 CP2_5_stage_0/charge_pump_1/capacitors_5_1/capacitor_5_3/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C892 CP2_5_stage_0/charge_pump_1/capacitors_5_1/capacitor_5_3/buffer_and_gate_0/in1 0 2.57f
C893 CP2_5_stage_0/charge_pump_1/capacitors_5_1/capacitor_5_2/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C894 CP2_5_stage_0/charge_pump_1/capacitors_5_1/capacitor_5_2/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C895 CP2_5_stage_0/charge_pump_1/capacitors_5_1/capacitor_5_2/buffer_and_gate_0/in1 0 2.57f
C896 CP2_5_stage_0/charge_pump_1/capacitors_5_1/capacitor_5_1/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C897 CP2_5_stage_0/charge_pump_1/capacitors_5_1/capacitor_5_1/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C898 CP2_5_stage_0/charge_pump_1/capacitors_5_1/capacitor_5_1/buffer_and_gate_0/in1 0 2.57f
C899 CP2_5_stage_0/charge_pump_1/capacitors_5_1/capacitor_5_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C900 CP2_5_stage_0/charge_pump_1/capacitors_5_1/capacitor_5_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C901 CP2_5_stage_0/charge_pump_1/capacitors_5_1/capacitor_5_0/buffer_and_gate_0/in1 0 2.57f
C902 CP2_5_stage_0/charge_pump_1/nmos_dnw3_0/out2 0 13.6f
C903 CP2_5_stage_0/charge_pump_1/capacitors_5_1/capacitor_5_7/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C904 CP2_5_stage_0/charge_pump_1/clock_0/clkb 0 80.5f
C905 CP2_5_stage_0/charge_pump_1/capacitors_5_1/capacitor_5_7/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C906 CP2_5_stage_0/charge_pump_1/capacitors_5_1/capacitor_5_7/buffer_and_gate_0/in1 0 2.57f
C907 CP2_5_stage_0/charge_pump_1/capacitors_5_1/capacitor_5_6/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C908 CP2_5_stage_0/charge_pump_1/capacitors_5_1/capacitor_5_6/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C909 CP2_5_stage_0/charge_pump_1/capacitors_5_1/capacitor_5_6/buffer_and_gate_0/in1 0 2.57f
C910 CP2_5_stage_0/charge_pump_1/capacitors_5_1/capacitor_5_5/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C911 CP2_5_stage_0/charge_pump_1/capacitors_5_1/capacitor_5_5/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C912 CP2_5_stage_0/charge_pump_1/capacitors_5_1/capacitor_5_5/buffer_and_gate_0/in1 0 2.57f
C913 CP2_5_stage_0/charge_pump_1/nmos_dnw3_0/clk 0 2.76f
C914 CP2_5_stage_0/charge_pump_0/nmos_dnw3_0/vs 0 16.4f
C915 CP2_5_stage_0/charge_pump_reverse_0/nmos_dnw3_0/vin 0 2.34f
C916 CP2_5_stage_0/charge_pump_0/clock_0/a_2432_n962# 0 8.68f **FLOATING
C917 CP2_5_stage_0/charge_pump_0/clock_0/a_2020_n482# 0 2.57f **FLOATING
C918 CP2_5_stage_0/charge_pump_0/clock_0/a_344_102# 0 2.81f
C919 CP2_5_stage_0/charge_pump_0/clock_0/a_2402_572# 0 2.17f
C920 CP2_5_stage_0/charge_pump_0/clock_0/a_344_n986# 0 2.38f
C921 CP2_5_stage_0/charge_pump_0/clock_0/clk_in 0 15.3f
C922 CP2_5_stage_0/charge_pump_0/clock_0/a_3246_118# 0 6.83f
C923 CP2_5_stage_0/charge_pump_0/nmos_dnw3_0/clkb 0 2.54f
C924 CP2_5_stage_0/charge_pump_0/capacitors_5_0/capacitor_5_4/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C925 CP2_5_stage_0/charge_pump_0/capacitors_5_0/capacitor_5_4/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C926 CP2_5_stage_0/charge_pump_0/capacitors_5_0/capacitor_5_4/buffer_and_gate_0/in1 0 2.57f
C927 CP2_5_stage_0/charge_pump_0/capacitors_5_0/capacitor_5_3/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C928 CP2_5_stage_0/charge_pump_0/capacitors_5_0/capacitor_5_3/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C929 CP2_5_stage_0/charge_pump_0/capacitors_5_0/capacitor_5_3/buffer_and_gate_0/in1 0 2.57f
C930 CP2_5_stage_0/charge_pump_0/capacitors_5_0/capacitor_5_2/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C931 CP2_5_stage_0/charge_pump_0/capacitors_5_0/capacitor_5_2/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C932 CP2_5_stage_0/charge_pump_0/capacitors_5_0/capacitor_5_2/buffer_and_gate_0/in1 0 2.57f
C933 CP2_5_stage_0/charge_pump_0/capacitors_5_0/capacitor_5_1/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C934 CP2_5_stage_0/charge_pump_0/capacitors_5_0/capacitor_5_1/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C935 CP2_5_stage_0/charge_pump_0/capacitors_5_0/capacitor_5_1/buffer_and_gate_0/in1 0 2.57f
C936 CP2_5_stage_0/charge_pump_0/capacitors_5_0/capacitor_5_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C937 CP2_5_stage_0/charge_pump_0/capacitors_5_0/capacitor_5_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C938 CP2_5_stage_0/charge_pump_0/capacitors_5_0/capacitor_5_0/buffer_and_gate_0/in1 0 2.57f
C939 CP2_5_stage_0/charge_pump_0/nmos_dnw3_0/out1 0 15f
C940 CP2_5_stage_0/charge_pump_0/capacitors_5_0/capacitor_5_7/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C941 CP2_5_stage_0/charge_pump_0/clock_0/clk 0 78.7f
C942 CP2_5_stage_0/charge_pump_0/capacitors_5_0/capacitor_5_7/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C943 CP2_5_stage_0/charge_pump_0/capacitors_5_0/capacitor_5_7/buffer_and_gate_0/in1 0 2.57f
C944 CP2_5_stage_0/charge_pump_0/capacitors_5_0/capacitor_5_6/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C945 CP2_5_stage_0/charge_pump_0/capacitors_5_0/capacitor_5_6/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C946 CP2_5_stage_0/charge_pump_0/capacitors_5_0/capacitor_5_6/buffer_and_gate_0/in1 0 2.57f
C947 scanchain_0/data_out[1] 0 23.6f
C948 CP2_5_stage_0/charge_pump_0/capacitors_5_0/capacitor_5_5/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C949 CP2_5_stage_0/charge_pump_0/capacitors_5_0/capacitor_5_5/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C950 CP2_5_stage_0/charge_pump_0/capacitors_5_0/capacitor_5_5/buffer_and_gate_0/in1 0 2.57f
C951 scanchain_0/data_out[2] 0 27.3f
C952 CP2_5_stage_0/charge_pump_0/capacitors_5_1/capacitor_5_4/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C953 CP2_5_stage_0/charge_pump_0/capacitors_5_1/capacitor_5_4/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C954 CP2_5_stage_0/charge_pump_0/capacitors_5_1/capacitor_5_4/buffer_and_gate_0/in1 0 2.57f
C955 CP2_5_stage_0/charge_pump_0/capacitors_5_1/capacitor_5_3/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C956 CP2_5_stage_0/charge_pump_0/capacitors_5_1/capacitor_5_3/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C957 CP2_5_stage_0/charge_pump_0/capacitors_5_1/capacitor_5_3/buffer_and_gate_0/in1 0 2.57f
C958 CP2_5_stage_0/charge_pump_0/capacitors_5_1/capacitor_5_2/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C959 CP2_5_stage_0/charge_pump_0/capacitors_5_1/capacitor_5_2/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C960 CP2_5_stage_0/charge_pump_0/capacitors_5_1/capacitor_5_2/buffer_and_gate_0/in1 0 2.57f
C961 CP2_5_stage_0/charge_pump_0/capacitors_5_1/capacitor_5_1/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C962 CP2_5_stage_0/charge_pump_0/capacitors_5_1/capacitor_5_1/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C963 CP2_5_stage_0/charge_pump_0/capacitors_5_1/capacitor_5_1/buffer_and_gate_0/in1 0 2.57f
C964 CP2_5_stage_0/charge_pump_0/capacitors_5_1/capacitor_5_0/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C965 CP2_5_stage_0/charge_pump_0/capacitors_5_1/capacitor_5_0/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C966 CP2_5_stage_0/charge_pump_0/capacitors_5_1/capacitor_5_0/buffer_and_gate_0/in1 0 2.57f
C967 CP2_5_stage_0/charge_pump_0/nmos_dnw3_0/out2 0 13.6f
C968 CP2_5_stage_0/charge_pump_0/capacitors_5_1/capacitor_5_7/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C969 CP2_5_stage_0/charge_pump_0/clock_0/clkb 0 80.5f
C970 CP2_5_stage_0/charge_pump_0/capacitors_5_1/capacitor_5_7/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C971 CP2_5_stage_0/charge_pump_0/capacitors_5_1/capacitor_5_7/buffer_and_gate_0/in1 0 2.57f
C972 CP2_5_stage_0/charge_pump_0/capacitors_5_1/capacitor_5_6/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C973 CP2_5_stage_0/charge_pump_0/capacitors_5_1/capacitor_5_6/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C974 CP2_5_stage_0/charge_pump_0/capacitors_5_1/capacitor_5_6/buffer_and_gate_0/in1 0 2.57f
C975 CP2_5_stage_0/charge_pump_0/capacitors_5_1/capacitor_5_5/buffer_and_gate_0/and_gate_0/a_n78_396# 0 2.34f
C976 CP2_5_stage_0/charge_pump_0/capacitors_5_1/capacitor_5_5/buffer_and_gate_0/buffer_0/a_1436_1552# 0 8.93f
C977 CP2_5_stage_0/charge_pump_0/capacitors_5_1/capacitor_5_5/buffer_and_gate_0/in1 0 2.57f
C978 CP2_5_stage_0/charge_pump_0/nmos_dnw3_0/clk 0 2.76f
.ends

