magic
tech sky130A
magscale 1 2
timestamp 1699074106
<< metal3 >>
rect -846 -14752 -624 894
rect 8778 734 9494 948
rect 9002 -14934 9494 734
<< metal4 >>
rect -1378 -14752 -806 1666
rect 7304 1474 9898 2028
rect 7448 -614 10042 -60
rect 7338 -2682 9932 -2128
rect 7434 -4776 10028 -4222
rect 7420 -6892 10014 -6338
rect 7462 -8946 10056 -8392
rect 7414 -11014 10008 -10460
rect 7462 -13116 10056 -12562
rect -1378 -14758 -1150 -14752
<< metal5 >>
rect -1972 -14744 -1314 569
rect 7420 2 10014 556
rect 7414 -2094 10008 -1540
rect 7358 -4168 9952 -3614
rect 7440 -6248 10034 -5694
rect 7414 -8330 10008 -7776
rect 7358 -10404 9952 -9850
rect 7420 -12520 10014 -11966
rect 7502 -14574 10096 -14020
use capacitor_5  capacitor_5_0
timestamp 1699074083
transform 1 0 0 0 1 18
box -1972 -346 8998 2050
use capacitor_5  capacitor_5_1
timestamp 1699074083
transform 1 0 12 0 1 -2068
box -1972 -346 8998 2050
use capacitor_5  capacitor_5_2
timestamp 1699074083
transform 1 0 14 0 1 -4162
box -1972 -346 8998 2050
use capacitor_5  capacitor_5_3
timestamp 1699074083
transform 1 0 88 0 1 -6252
box -1972 -346 8998 2050
use capacitor_5  capacitor_5_4
timestamp 1699074083
transform 1 0 88 0 1 -8350
box -1972 -346 8998 2050
use capacitor_5  capacitor_5_5
timestamp 1699074083
transform 1 0 88 0 1 -10432
box -1972 -346 8998 2050
use capacitor_5  capacitor_5_6
timestamp 1699074083
transform 1 0 86 0 1 -12526
box -1972 -346 8998 2050
use capacitor_5  capacitor_5_7
timestamp 1699074083
transform 1 0 86 0 1 -14612
box -1972 -346 8998 2050
<< end >>
