magic
tech sky130A
magscale 1 2
timestamp 1698389451
<< nwell >>
rect 610 760 862 762
rect 564 758 1076 760
rect 564 754 1556 758
rect -260 290 1556 754
rect -260 286 1348 290
<< nmos >>
rect -16 -64 14 20
rect 80 -64 110 20
rect 176 -64 206 20
rect 272 -64 302 20
rect 368 -64 398 20
rect 464 -64 494 20
rect 556 -64 586 20
<< pmos >>
rect -16 396 14 648
rect 80 396 110 648
rect 176 396 206 648
rect 272 396 302 648
rect 368 396 398 648
rect 464 396 494 648
rect 556 396 586 648
<< ndiff >>
rect -78 8 -16 20
rect -78 -52 -66 8
rect -32 -52 -16 8
rect -78 -64 -16 -52
rect 14 8 80 20
rect 14 -52 30 8
rect 64 -52 80 8
rect 14 -64 80 -52
rect 110 8 176 20
rect 110 -52 126 8
rect 160 -52 176 8
rect 110 -64 176 -52
rect 206 8 272 20
rect 206 -52 222 8
rect 256 -52 272 8
rect 206 -64 272 -52
rect 302 8 368 20
rect 302 -52 318 8
rect 352 -52 368 8
rect 302 -64 368 -52
rect 398 8 464 20
rect 398 -52 414 8
rect 448 -52 464 8
rect 398 -64 464 -52
rect 494 8 556 20
rect 494 -52 510 8
rect 544 -52 556 8
rect 494 -64 556 -52
rect 586 8 644 20
rect 586 -52 598 8
rect 632 -52 644 8
rect 586 -64 644 -52
<< pdiff >>
rect -78 636 -16 648
rect -78 408 -66 636
rect -32 408 -16 636
rect -78 396 -16 408
rect 14 636 80 648
rect 14 408 30 636
rect 64 408 80 636
rect 14 396 80 408
rect 110 636 176 648
rect 110 408 126 636
rect 160 408 176 636
rect 110 396 176 408
rect 206 636 272 648
rect 206 408 222 636
rect 256 408 272 636
rect 206 396 272 408
rect 302 636 368 648
rect 302 408 318 636
rect 352 408 368 636
rect 302 396 368 408
rect 398 636 464 648
rect 398 408 414 636
rect 448 408 464 636
rect 398 396 464 408
rect 494 636 556 648
rect 494 408 510 636
rect 544 408 556 636
rect 494 396 556 408
rect 586 636 644 648
rect 586 408 598 636
rect 632 408 644 636
rect 586 396 644 408
<< ndiffc >>
rect -66 -52 -32 8
rect 30 -52 64 8
rect 126 -52 160 8
rect 222 -52 256 8
rect 318 -52 352 8
rect 414 -52 448 8
rect 510 -52 544 8
rect 598 -52 632 8
<< pdiffc >>
rect -66 408 -32 636
rect 30 408 64 636
rect 126 408 160 636
rect 222 408 256 636
rect 318 408 352 636
rect 414 408 448 636
rect 510 408 544 636
rect 598 408 632 636
<< psubdiff >>
rect -220 6 -132 20
rect -220 -50 -194 6
rect -156 -50 -132 6
rect -220 -64 -132 -50
<< nsubdiff >>
rect -224 628 -142 654
rect -224 414 -200 628
rect -166 414 -142 628
rect -224 384 -142 414
<< psubdiffcont >>
rect -194 -50 -156 6
<< nsubdiffcont >>
rect -200 414 -166 628
<< poly >>
rect -34 729 32 745
rect -34 695 -18 729
rect 16 728 32 729
rect 158 729 224 745
rect 158 728 174 729
rect 16 695 174 728
rect 208 728 224 729
rect 350 729 416 745
rect 350 728 366 729
rect 208 695 366 728
rect 400 728 416 729
rect 400 695 496 728
rect -34 694 496 695
rect 798 696 1328 730
rect -34 679 32 694
rect -16 648 14 679
rect 80 648 110 694
rect 158 679 224 694
rect 176 648 206 679
rect 272 648 302 694
rect 350 679 416 694
rect 368 648 398 679
rect 464 648 494 694
rect 556 648 586 674
rect 798 652 828 696
rect 990 656 1020 696
rect 1182 650 1212 696
rect -16 352 14 396
rect 80 366 110 396
rect -24 348 14 352
rect 56 349 128 366
rect 176 354 206 396
rect 272 365 302 396
rect 254 364 320 365
rect 56 348 74 349
rect -24 315 74 348
rect 108 348 128 349
rect 172 348 206 354
rect 250 349 320 364
rect 250 348 266 349
rect 108 315 266 348
rect 300 348 320 349
rect 368 348 398 396
rect 464 366 494 396
rect 442 349 512 366
rect 442 348 458 349
rect 300 315 458 348
rect 492 315 512 349
rect -24 314 512 315
rect -24 266 10 314
rect 58 299 124 314
rect 250 299 316 314
rect 442 298 512 314
rect -162 254 10 266
rect -162 216 -146 254
rect -6 218 10 254
rect -6 216 12 218
rect -162 206 12 216
rect -24 108 12 206
rect 556 200 586 396
rect 794 348 828 352
rect 894 348 924 390
rect 1086 348 1116 388
rect 1278 348 1308 388
rect 780 314 1308 348
rect 794 238 828 314
rect 634 226 828 238
rect 514 184 588 200
rect 514 150 538 184
rect 572 150 588 184
rect 634 188 650 226
rect 812 188 828 226
rect 634 178 828 188
rect 514 134 588 150
rect -34 92 32 108
rect 158 92 224 108
rect 350 92 416 108
rect -34 58 -18 92
rect 16 58 174 92
rect 208 58 366 92
rect 400 58 494 92
rect -34 42 32 58
rect -16 20 14 42
rect 80 20 110 58
rect 158 42 224 58
rect 176 20 206 42
rect 272 20 302 58
rect 350 42 416 58
rect 368 20 398 42
rect 464 20 494 58
rect 556 20 586 134
rect 794 100 828 178
rect 794 70 1326 100
rect 798 62 1326 70
rect 798 30 828 62
rect 990 40 1020 62
rect 1182 40 1212 62
rect -16 -102 14 -64
rect 80 -86 110 -64
rect 62 -102 128 -86
rect 176 -102 206 -64
rect 272 -86 302 -64
rect 254 -102 320 -86
rect 368 -102 398 -64
rect 464 -86 494 -64
rect 446 -102 512 -86
rect 556 -90 586 -64
rect 894 -98 924 -68
rect 1086 -98 1116 -68
rect 1278 -98 1308 -64
rect -16 -134 78 -102
rect 62 -136 78 -134
rect 112 -134 270 -102
rect 112 -136 128 -134
rect 62 -152 128 -136
rect 254 -136 270 -134
rect 304 -134 462 -102
rect 304 -136 320 -134
rect 254 -152 320 -136
rect 446 -136 462 -134
rect 496 -136 512 -102
rect 780 -132 1308 -98
rect 446 -152 512 -136
<< polycont >>
rect -18 695 16 729
rect 174 695 208 729
rect 366 695 400 729
rect 74 315 108 349
rect 266 315 300 349
rect 458 315 492 349
rect -146 216 -6 254
rect 538 150 572 184
rect 650 188 812 226
rect -18 58 16 92
rect 174 58 208 92
rect 366 58 400 92
rect 78 -136 112 -102
rect 270 -136 304 -102
rect 462 -136 496 -102
<< locali >>
rect -34 695 -18 729
rect 16 695 32 729
rect 158 695 174 729
rect 208 695 224 729
rect 350 695 366 729
rect 400 695 416 729
rect -216 628 -150 646
rect -216 414 -200 628
rect -166 414 -150 628
rect -216 394 -150 414
rect -66 636 -32 652
rect -66 392 -32 408
rect 30 636 64 652
rect 30 392 64 408
rect 126 636 160 652
rect 126 392 160 408
rect 222 636 256 652
rect 222 392 256 408
rect 318 636 352 652
rect 318 392 352 408
rect 414 636 448 652
rect 414 392 448 408
rect 510 636 544 652
rect 510 392 544 408
rect 598 636 632 652
rect 598 392 632 408
rect 58 315 74 349
rect 108 315 124 349
rect 250 315 266 349
rect 300 315 316 349
rect 442 315 458 349
rect 492 315 508 349
rect -260 268 12 282
rect -260 216 -246 268
rect -62 266 12 268
rect -8 254 12 266
rect -6 216 12 254
rect -260 208 12 216
rect -164 204 12 208
rect 634 226 828 238
rect 404 184 590 200
rect 404 148 428 184
rect 572 148 590 184
rect 634 188 650 226
rect 812 188 828 226
rect 634 178 828 188
rect 404 134 590 148
rect -34 58 -18 92
rect 16 58 32 92
rect 158 58 174 92
rect 208 58 224 92
rect 350 58 366 92
rect 400 58 416 92
rect -66 12 -32 24
rect -214 6 -132 12
rect -214 -50 -194 6
rect -156 -50 -132 6
rect -214 -56 -132 -50
rect -78 8 -32 12
rect -78 -52 -66 8
rect -78 -56 -32 -52
rect -66 -68 -32 -56
rect 30 8 64 24
rect 30 -68 64 -52
rect 126 8 160 24
rect 126 -68 160 -52
rect 222 8 256 24
rect 222 -68 256 -52
rect 318 8 352 24
rect 318 -68 352 -52
rect 414 8 448 24
rect 414 -68 448 -52
rect 510 8 544 24
rect 510 -68 544 -52
rect 598 8 632 24
rect 598 -68 632 -52
rect 62 -136 78 -102
rect 112 -136 128 -102
rect 254 -136 270 -102
rect 304 -136 320 -102
rect 446 -136 462 -102
rect 496 -136 512 -102
<< viali >>
rect -200 414 -166 628
rect -66 408 -32 636
rect 30 408 64 636
rect 126 408 160 636
rect 222 408 256 636
rect 318 408 352 636
rect 414 408 448 636
rect 510 408 544 636
rect 598 408 632 636
rect -246 266 -62 268
rect -246 254 -8 266
rect -246 216 -146 254
rect -146 216 -6 254
rect 428 150 538 184
rect 538 150 572 184
rect 428 148 572 150
rect 650 188 812 226
rect -194 -50 -156 6
rect -66 -52 -32 8
rect 30 -52 64 8
rect 126 -52 160 8
rect 222 -52 256 8
rect 318 -52 352 8
rect 414 -52 448 8
rect 510 -52 544 8
rect 598 -52 632 8
<< metal1 >>
rect -684 1272 1674 1316
rect -684 804 -620 1272
rect 1594 1254 1674 1272
rect -684 786 -614 804
rect 1600 786 1674 1254
rect -684 772 1674 786
rect -216 770 1260 772
rect -216 768 876 770
rect -216 760 634 768
rect -216 628 -150 760
rect -86 648 -16 652
rect 28 648 64 760
rect -216 414 -200 628
rect -166 414 -150 628
rect -216 396 -150 414
rect -88 638 -16 648
rect -88 408 -78 638
rect -18 408 -16 638
rect -88 404 -16 408
rect 24 636 70 648
rect 24 408 30 636
rect 64 408 70 636
rect -88 400 -18 404
rect -72 396 -26 400
rect 24 396 70 408
rect 106 638 176 650
rect 222 648 258 760
rect 414 648 450 760
rect 106 408 112 638
rect 172 408 176 638
rect 106 402 176 408
rect 216 636 262 648
rect 216 408 222 636
rect 256 408 262 636
rect 120 396 166 402
rect 216 396 262 408
rect 300 638 370 648
rect 300 408 308 638
rect 368 408 370 638
rect 300 400 370 408
rect 408 636 454 648
rect 408 408 414 636
rect 448 408 454 636
rect 312 396 358 400
rect 408 396 454 408
rect 494 636 564 650
rect 598 648 634 760
rect 494 410 500 636
rect 556 410 564 636
rect 494 408 510 410
rect 544 408 564 410
rect 494 402 564 408
rect 592 636 638 648
rect 592 408 598 636
rect 632 408 638 636
rect 844 514 876 768
rect 1038 518 1070 770
rect 1228 514 1260 770
rect 504 396 550 402
rect 592 396 638 408
rect -68 394 -34 396
rect 124 394 158 396
rect 318 394 352 396
rect 510 394 544 396
rect 748 362 782 424
rect 940 362 974 428
rect 748 328 974 362
rect -260 268 12 282
rect -260 216 -246 268
rect 6 216 12 268
rect -260 214 -146 216
rect -6 214 12 216
rect -260 208 12 214
rect 622 236 828 238
rect 404 184 590 200
rect 404 178 428 184
rect -134 148 428 178
rect 572 148 590 184
rect 622 184 650 236
rect 812 184 828 236
rect 622 178 828 184
rect 940 150 974 328
rect 1132 150 1166 424
rect 1324 150 1358 430
rect -132 134 590 148
rect 748 118 1360 150
rect -86 20 -16 26
rect -212 6 -138 12
rect -212 -50 -194 6
rect -156 -50 -138 6
rect -212 -56 -138 -50
rect -203 -156 -169 -56
rect -86 -64 -78 20
rect -22 -64 -16 20
rect 24 8 70 20
rect 24 -52 30 8
rect 64 -52 70 8
rect 24 -64 70 -52
rect 108 10 178 26
rect 316 24 350 26
rect 510 24 544 26
rect 108 -52 116 10
rect 168 -52 178 10
rect -86 -66 -16 -64
rect 30 -156 64 -64
rect 108 -66 178 -52
rect 216 8 262 20
rect 216 -52 222 8
rect 256 -52 262 8
rect 216 -64 262 -52
rect 302 8 372 24
rect 302 -54 308 8
rect 360 -54 372 8
rect -203 -158 64 -156
rect 222 -158 256 -64
rect 302 -68 372 -54
rect 408 8 454 20
rect 408 -52 414 8
rect 448 -52 454 8
rect 408 -64 454 -52
rect 494 8 556 24
rect 592 18 642 20
rect 494 -54 500 8
rect 552 -54 556 8
rect 414 -158 448 -64
rect 494 -66 556 -54
rect 584 8 644 18
rect 584 -54 588 8
rect 642 -54 644 8
rect 748 -50 782 118
rect 584 -62 644 -54
rect 592 -64 638 -62
rect 844 -158 878 10
rect 940 -50 974 118
rect 1036 -158 1070 10
rect 1132 -50 1166 118
rect 1228 -158 1262 10
rect 1324 -50 1358 118
rect -204 -166 1262 -158
rect -204 -230 -192 -166
rect 1252 -230 1262 -166
rect -204 -246 1262 -230
<< via1 >>
rect -620 1254 1594 1272
rect -620 804 1600 1254
rect -614 786 1600 804
rect -78 636 -18 638
rect -78 408 -66 636
rect -66 408 -32 636
rect -32 408 -18 636
rect 112 636 172 638
rect 112 408 126 636
rect 126 408 160 636
rect 160 408 172 636
rect 308 636 368 638
rect 308 408 318 636
rect 318 408 352 636
rect 352 408 368 636
rect 500 410 510 636
rect 510 410 544 636
rect 544 410 556 636
rect -246 266 -62 268
rect -62 266 6 268
rect -246 254 -8 266
rect -8 254 6 266
rect -246 216 -6 254
rect -6 216 6 254
rect -146 214 -6 216
rect 650 226 812 236
rect 650 188 812 226
rect 650 184 812 188
rect -78 8 -22 20
rect -78 -52 -66 8
rect -66 -52 -32 8
rect -32 -52 -22 8
rect -78 -64 -22 -52
rect 116 8 168 10
rect 116 -52 126 8
rect 126 -52 160 8
rect 160 -52 168 8
rect 308 -52 318 8
rect 318 -52 352 8
rect 352 -52 360 8
rect 308 -54 360 -52
rect 500 -52 510 8
rect 510 -52 544 8
rect 544 -52 552 8
rect 500 -54 552 -52
rect 588 -52 598 8
rect 598 -52 632 8
rect 632 -52 642 8
rect 588 -54 642 -52
rect -192 -230 1252 -166
<< metal2 >>
rect -684 1272 1674 1316
rect -684 804 -620 1272
rect 1594 1254 1674 1272
rect -684 786 -614 804
rect 1600 786 1674 1254
rect -684 772 1674 786
rect -88 638 566 650
rect -88 408 -78 638
rect -18 408 112 638
rect 172 408 308 638
rect 368 636 566 638
rect 368 408 496 636
rect 560 408 566 636
rect -88 402 566 408
rect 486 398 566 402
rect 508 392 546 398
rect -256 282 -216 286
rect -260 280 -162 282
rect -122 280 12 282
rect -260 268 12 280
rect -260 216 -246 268
rect 6 216 12 268
rect -260 214 -146 216
rect -6 214 12 216
rect -260 204 12 214
rect 634 236 828 238
rect 634 180 650 236
rect 812 180 828 236
rect 634 178 828 180
rect -86 20 554 22
rect -86 -64 -78 20
rect -22 10 554 20
rect -22 -52 116 10
rect 168 8 554 10
rect 168 -52 308 8
rect -22 -54 308 -52
rect 360 -54 500 8
rect 552 -54 554 8
rect -22 -64 554 -54
rect 584 8 646 26
rect 584 -54 588 8
rect 644 -54 646 8
rect 584 -64 646 -54
rect -204 -164 1262 -158
rect -204 -230 -192 -164
rect 1252 -230 1262 -164
rect -204 -246 1262 -230
<< via2 >>
rect -620 1254 1594 1272
rect -620 804 1600 1254
rect -614 786 1600 804
rect 496 410 500 636
rect 500 410 556 636
rect 556 410 560 636
rect 496 408 560 410
rect 650 184 812 236
rect 650 180 812 184
rect 588 -54 642 8
rect 642 -54 644 8
rect -192 -166 1252 -164
rect -192 -230 1252 -166
<< metal3 >>
rect -684 1272 1674 1316
rect -684 804 -620 1272
rect 1594 1254 1674 1272
rect -684 786 -614 804
rect 1600 786 1674 1254
rect -684 772 1674 786
rect 486 636 566 650
rect 486 408 496 636
rect 560 408 566 636
rect 486 398 566 408
rect 496 268 562 398
rect 496 242 644 268
rect 496 236 828 242
rect 496 196 650 236
rect 584 180 650 196
rect 812 180 828 236
rect 584 172 828 180
rect 584 26 644 172
rect 578 8 652 26
rect 578 -54 588 8
rect 644 -54 652 8
rect 578 -62 652 -54
rect 584 -64 646 -62
rect -204 -164 1262 -158
rect -204 -230 -192 -164
rect 1252 -230 1262 -164
rect -204 -246 1262 -230
<< via3 >>
rect -620 1254 1594 1272
rect -620 804 1600 1254
rect -614 786 1600 804
rect -192 -230 1252 -166
<< metal4 >>
rect -684 1272 1674 1316
rect -684 804 -620 1272
rect 1594 1254 1674 1272
rect -684 786 -614 804
rect 1600 786 1674 1254
rect -684 772 1674 786
rect -676 -166 1688 -150
rect -676 -230 -192 -166
rect 1252 -230 1688 -166
rect -676 -258 1688 -230
rect -676 -598 -552 -258
rect 1566 -598 1688 -258
rect -676 -688 1688 -598
<< via4 >>
rect -552 -598 1566 -258
<< metal5 >>
rect -676 -258 1688 -150
rect -676 -598 -552 -258
rect 1566 -598 1688 -258
rect -676 -688 1688 -598
use sky130_fd_pr__nfet_01v8_XJUN3E  sky130_fd_pr__nfet_01v8_XJUN3E_0 ~/Desktop/charge_pumps2/layout_files
timestamp 1697701953
transform 1 0 1053 0 1 -20
box -317 -130 317 130
use sky130_fd_pr__pfet_01v8_X4L24Q  sky130_fd_pr__pfet_01v8_X4L24Q_0 ~/Desktop/charge_pumps2/layout_files
timestamp 1697701953
transform 1 0 1053 0 1 522
box -353 -226 353 226
<< end >>
