magic
tech sky130A
magscale 1 2
timestamp 1698760865
<< nwell >>
rect 20588 -2182 21342 -1808
rect 26126 -2168 26790 -1790
rect 45066 -2094 45282 -1720
rect 47354 -2104 47944 -1728
rect 68172 -2050 68860 -1674
rect 70956 -2036 71258 -1660
rect 91412 -2132 91748 -1756
rect 93910 -2110 94136 -1734
<< nsubdiff >>
rect 68662 -1870 68762 -1840
rect 21112 -1952 21228 -1914
rect 21112 -2042 21138 -1952
rect 21194 -2042 21228 -1952
rect 45122 -1918 45208 -1888
rect 45122 -1960 45148 -1918
rect 45186 -1960 45208 -1918
rect 21112 -2100 21228 -2042
rect 26216 -1988 26308 -1962
rect 45122 -1984 45208 -1960
rect 47390 -1904 47484 -1876
rect 47390 -1944 47418 -1904
rect 47454 -1944 47484 -1904
rect 68662 -1906 68686 -1870
rect 68728 -1906 68762 -1870
rect 68662 -1930 68762 -1906
rect 71022 -1846 71116 -1824
rect 71022 -1886 71048 -1846
rect 71090 -1886 71116 -1846
rect 71022 -1910 71116 -1886
rect 91522 -1926 91630 -1900
rect 47390 -1968 47484 -1944
rect 91522 -1968 91548 -1926
rect 91604 -1968 91630 -1926
rect 26216 -2022 26244 -1988
rect 26280 -2022 26308 -1988
rect 91522 -1994 91630 -1968
rect 93976 -1918 94072 -1892
rect 93976 -1964 93998 -1918
rect 94040 -1964 94072 -1918
rect 93976 -1990 94072 -1964
rect 26216 -2048 26308 -2022
<< nsubdiffcont >>
rect 21138 -2042 21194 -1952
rect 45148 -1960 45186 -1918
rect 47418 -1944 47454 -1904
rect 68686 -1906 68728 -1870
rect 71048 -1886 71090 -1846
rect 91548 -1968 91604 -1926
rect 26244 -2022 26280 -1988
rect 93998 -1964 94040 -1918
<< locali >>
rect 68662 -1870 68762 -1840
rect 21112 -1952 21228 -1914
rect 21112 -2042 21138 -1952
rect 21194 -2042 21228 -1952
rect 45122 -1918 45208 -1888
rect 45122 -1960 45148 -1918
rect 45186 -1960 45208 -1918
rect 21112 -2100 21228 -2042
rect 26216 -1988 26308 -1962
rect 45122 -1984 45208 -1960
rect 47390 -1904 47484 -1876
rect 47390 -1944 47418 -1904
rect 47454 -1944 47484 -1904
rect 68662 -1906 68686 -1870
rect 68728 -1906 68762 -1870
rect 68662 -1930 68762 -1906
rect 71022 -1846 71116 -1824
rect 71022 -1886 71048 -1846
rect 71090 -1886 71116 -1846
rect 71022 -1910 71116 -1886
rect 91522 -1926 91630 -1900
rect 47390 -1968 47484 -1944
rect 91522 -1968 91548 -1926
rect 91604 -1968 91630 -1926
rect 26216 -2022 26244 -1988
rect 26280 -2022 26308 -1988
rect 91522 -1994 91630 -1968
rect 93976 -1918 94072 -1892
rect 93976 -1964 93998 -1918
rect 94040 -1964 94072 -1918
rect 93976 -1990 94072 -1964
rect 26216 -2048 26308 -2022
<< viali >>
rect 21138 -2042 21194 -1952
rect 45148 -1960 45186 -1918
rect 47418 -1944 47454 -1904
rect 68686 -1906 68728 -1870
rect 71048 -1886 71090 -1846
rect 91548 -1968 91604 -1926
rect 26244 -2022 26280 -1988
rect 93998 -1964 94040 -1918
<< metal1 >>
rect 19362 -1277 26746 -1232
rect 19350 -1823 26761 -1277
rect 43315 -1726 47861 -1443
rect 66304 -1670 71488 -1470
rect 26990 -1818 27382 -1766
rect 19350 -2622 19896 -1823
rect 21138 -1914 21196 -1823
rect 21112 -1952 21228 -1914
rect 21112 -2042 21138 -1952
rect 21194 -2042 21228 -1952
rect 26244 -1962 26282 -1823
rect 21112 -2100 21228 -2042
rect 26216 -1988 26308 -1962
rect 26216 -2022 26244 -1988
rect 26280 -2022 26308 -1988
rect 26216 -2048 26308 -2022
rect 20940 -2176 26150 -2150
rect 26990 -2169 27042 -1818
rect 20940 -2204 26166 -2176
rect 26708 -2203 27042 -2169
rect 20940 -2218 26150 -2204
rect 21010 -2222 26150 -2218
rect 26990 -2268 27042 -2203
rect 27336 -2268 27382 -1818
rect 26990 -2316 27382 -2268
rect 20634 -2376 20668 -2324
rect 20852 -2376 20886 -2324
rect 26402 -2376 26436 -2336
rect 26620 -2376 26654 -2336
rect 26945 -2376 27138 -2372
rect 19004 -2722 20346 -2622
rect 19004 -3184 19172 -2722
rect 20150 -3184 20346 -2722
rect 20606 -2922 27138 -2376
rect 43315 -2606 43437 -1726
rect 45148 -1888 45186 -1726
rect 47418 -1876 47456 -1726
rect 47982 -1830 48384 -1758
rect 45122 -1918 45208 -1888
rect 45122 -1960 45148 -1918
rect 45186 -1960 45208 -1918
rect 45122 -1984 45208 -1960
rect 47390 -1904 47484 -1876
rect 47390 -1944 47418 -1904
rect 47454 -1944 47484 -1904
rect 47390 -1968 47484 -1944
rect 45014 -2098 47370 -2094
rect 45044 -2122 47370 -2098
rect 47982 -2104 48050 -1830
rect 47926 -2106 48050 -2104
rect 47884 -2139 48050 -2106
rect 47982 -2172 48050 -2139
rect 48308 -2172 48384 -1830
rect 47982 -2224 48384 -2172
rect 44678 -2298 44712 -2242
rect 44896 -2298 44930 -2242
rect 47554 -2298 47588 -2252
rect 47772 -2298 47806 -2252
rect 44678 -2463 51541 -2298
rect 44686 -2464 51541 -2463
rect 19004 -3278 20346 -3184
rect 26592 -3868 27138 -2922
rect 42944 -2686 44082 -2606
rect 42944 -3226 43016 -2686
rect 43986 -3226 44082 -2686
rect 42944 -3268 44082 -3226
rect 43315 -3273 43437 -3268
rect 26394 -3990 27668 -3868
rect 51375 -3874 51541 -2464
rect 66304 -2618 66504 -1670
rect 68686 -1840 68730 -1670
rect 71048 -1824 71090 -1670
rect 89760 -1754 94436 -1586
rect 68662 -1870 68762 -1840
rect 68662 -1906 68686 -1870
rect 68728 -1906 68762 -1870
rect 68662 -1930 68762 -1906
rect 71022 -1846 71116 -1824
rect 71022 -1886 71048 -1846
rect 71090 -1886 71116 -1846
rect 71022 -1910 71116 -1886
rect 71622 -1830 72018 -1762
rect 71622 -2034 71670 -1830
rect 68586 -2076 71064 -2048
rect 71529 -2069 71670 -2034
rect 71622 -2146 71670 -2069
rect 71936 -2146 72018 -1830
rect 68216 -2272 68250 -2196
rect 71622 -2218 72018 -2146
rect 74451 -2272 74648 -2264
rect 68216 -2419 74651 -2272
rect 65758 -2732 67080 -2618
rect 65758 -3166 65848 -2732
rect 66898 -3166 67080 -2732
rect 65758 -3258 67080 -3166
rect 66378 -3288 66494 -3258
rect 26394 -4446 26522 -3990
rect 27568 -4446 27668 -3990
rect 26394 -4526 27668 -4446
rect 50940 -3928 51898 -3874
rect 74451 -3886 74648 -2419
rect 89760 -2626 89928 -1754
rect 91548 -1900 91604 -1754
rect 93998 -1892 94042 -1754
rect 94588 -1804 94996 -1754
rect 91522 -1926 91630 -1900
rect 91522 -1968 91548 -1926
rect 91604 -1968 91630 -1926
rect 91522 -1994 91630 -1968
rect 93976 -1918 94072 -1892
rect 93976 -1964 93998 -1918
rect 94040 -1964 94072 -1918
rect 93976 -1990 94072 -1964
rect 94588 -2108 94660 -1804
rect 91387 -2158 94078 -2130
rect 94493 -2143 94660 -2108
rect 91387 -2165 91491 -2158
rect 94588 -2230 94660 -2143
rect 94952 -2230 94996 -1804
rect 91074 -2324 91108 -2278
rect 91292 -2324 91326 -2278
rect 94164 -2324 94198 -2256
rect 94382 -2324 94416 -2256
rect 94588 -2284 94996 -2230
rect 91074 -2465 98420 -2324
rect 90368 -2626 90536 -2612
rect 89696 -2722 91328 -2626
rect 89696 -3208 89834 -2722
rect 91108 -3208 91328 -2722
rect 89696 -3304 91328 -3208
rect 90471 -3334 90505 -3304
rect 98279 -3886 98420 -2465
rect 50940 -4472 51026 -3928
rect 51844 -4472 51898 -3928
rect 50940 -4526 51898 -4472
rect 73315 -4010 75340 -3886
rect 73315 -4448 73494 -4010
rect 75202 -4448 75340 -4010
rect 73315 -4529 75340 -4448
rect 97388 -4008 99380 -3886
rect 97388 -4410 97540 -4008
rect 99214 -4410 99380 -4008
rect 97388 -4522 99380 -4410
rect 98341 -4527 98375 -4522
rect 74451 -4546 74648 -4529
<< via1 >>
rect 27042 -2268 27336 -1818
rect 19172 -3184 20150 -2722
rect 48050 -2172 48308 -1830
rect 43016 -3226 43986 -2686
rect 71670 -2146 71936 -1830
rect 65848 -3166 66898 -2732
rect 26522 -4446 27568 -3990
rect 94660 -2230 94952 -1804
rect 89834 -3208 91108 -2722
rect 51026 -4472 51844 -3928
rect 73494 -4448 75202 -4010
rect 97540 -4410 99214 -4008
<< metal2 >>
rect 44480 25420 46872 25660
rect 46632 24910 46872 25420
rect 91012 25410 94204 25650
rect 93964 24900 94204 25410
rect 25044 23722 25284 23734
rect 21716 23660 25284 23722
rect 45020 23670 48556 23726
rect 68452 23672 71968 23732
rect 25044 23594 25284 23660
rect 91694 23658 95834 23720
rect 21738 21584 25270 21646
rect 45036 21578 48572 21634
rect 68438 21574 71954 21634
rect 91682 21576 95822 21638
rect 21710 19618 21884 19626
rect 21710 19566 21916 19618
rect 21710 19510 25350 19566
rect 21728 19482 25350 19510
rect 45028 19492 48564 19548
rect 68426 19482 71942 19542
rect 91690 19482 95830 19544
rect 21636 17470 21828 17502
rect 21636 17442 25294 17470
rect 21636 17386 25328 17442
rect 45018 17406 48554 17462
rect 68360 17400 71876 17460
rect 91690 17386 95830 17448
rect 25056 17328 25328 17386
rect 21662 15314 25284 15398
rect 45020 15304 48556 15360
rect 68350 15302 71866 15362
rect 91686 15288 95826 15350
rect 21636 13224 25186 13270
rect 45102 13208 48610 13278
rect 68358 13218 71874 13278
rect 91774 13212 95914 13274
rect 21742 11118 25124 11190
rect 45096 11114 48604 11184
rect 68358 11120 71874 11180
rect 91760 11118 95900 11180
rect 21678 9032 25060 9104
rect 45096 9026 48604 9096
rect 68358 9026 71854 9106
rect 91764 9020 95904 9082
rect 23392 7344 23572 7974
rect 69950 7346 70190 7952
rect 11784 7104 23578 7344
rect 67368 7106 70190 7346
rect 26990 -1818 27382 -1766
rect 20148 -1950 20550 -1888
rect 20148 -2262 20198 -1950
rect 20512 -2150 20550 -1950
rect 20512 -2228 20574 -2150
rect 20512 -2262 20550 -2228
rect 20148 -2312 20550 -2262
rect 26990 -2268 27042 -1818
rect 27336 -2268 27382 -1818
rect 26990 -2316 27382 -2268
rect 43858 -1826 44494 -1754
rect 43858 -2250 43934 -1826
rect 44408 -2250 44494 -1826
rect 47982 -1830 48384 -1758
rect 47982 -2172 48050 -1830
rect 48308 -2172 48384 -1830
rect 47982 -2224 48384 -2172
rect 67564 -1786 68060 -1752
rect 43858 -2318 44494 -2250
rect 67564 -2272 67596 -1786
rect 68018 -2272 68060 -1786
rect 71622 -1830 72018 -1762
rect 94592 -1804 95002 -1754
rect 71622 -2146 71670 -1830
rect 71936 -2146 72018 -1830
rect 71622 -2218 72018 -2146
rect 90468 -1876 91004 -1818
rect 67564 -2316 68060 -2272
rect 90468 -2244 90546 -1876
rect 90922 -2244 91004 -1876
rect 90468 -2298 91004 -2244
rect 94592 -2230 94660 -1804
rect 94952 -2230 95002 -1804
rect 94592 -2290 95002 -2230
rect 19004 -2722 20346 -2622
rect 19004 -3184 19172 -2722
rect 20150 -3184 20346 -2722
rect 19004 -3278 20346 -3184
rect 42944 -2686 44082 -2606
rect 42944 -3226 43016 -2686
rect 43986 -3226 44082 -2686
rect 42944 -3268 44082 -3226
rect 65758 -2732 67080 -2618
rect 65758 -3166 65848 -2732
rect 66898 -3166 67080 -2732
rect 65758 -3258 67080 -3166
rect 89696 -2722 91328 -2626
rect 89696 -3208 89834 -2722
rect 91108 -3208 91328 -2722
rect 89696 -3304 91328 -3208
rect 26394 -3990 27668 -3868
rect 26394 -4446 26522 -3990
rect 27568 -4446 27668 -3990
rect 26394 -4526 27668 -4446
rect 50940 -3928 51898 -3874
rect 50940 -4472 51026 -3928
rect 51844 -4472 51898 -3928
rect 50940 -4526 51898 -4472
rect 73315 -4010 75340 -3886
rect 73315 -4448 73494 -4010
rect 75202 -4448 75340 -4010
rect 73315 -4529 75340 -4448
rect 97388 -4008 99380 -3886
rect 97388 -4410 97540 -4008
rect 99214 -4410 99380 -4008
rect 97388 -4522 99380 -4410
<< via2 >>
rect 20198 -2262 20512 -1950
rect 27042 -2268 27336 -1818
rect 43934 -2250 44408 -1826
rect 48050 -2172 48308 -1830
rect 67596 -2272 68018 -1786
rect 71670 -2146 71936 -1830
rect 90546 -2244 90922 -1876
rect 94660 -2230 94952 -1804
rect 19172 -3184 20150 -2722
rect 43016 -3226 43986 -2686
rect 65848 -3166 66898 -2732
rect 89834 -3208 91108 -2722
rect 26522 -4446 27568 -3990
rect 51026 -4472 51844 -3928
rect 73494 -4448 75202 -4010
rect 97540 -4410 99214 -4008
<< metal3 >>
rect 11892 -1760 11964 294
rect 17014 -1760 17084 -1756
rect 34918 -1760 34990 -766
rect 58636 -1760 58708 296
rect 67212 -1760 67278 -1738
rect 74954 -1760 75026 -1738
rect 94592 -1760 95002 -1754
rect -2079 -1950 20673 -1760
rect 26990 -1768 27382 -1766
rect 29650 -1768 44587 -1760
rect -2079 -2262 20198 -1950
rect 20512 -2262 20673 -1950
rect -2079 -2314 20673 -2262
rect 26779 -1818 44587 -1768
rect 26779 -2268 27042 -1818
rect 27336 -1826 44587 -1818
rect 27336 -2250 43934 -1826
rect 44408 -2250 44587 -1826
rect 27336 -2268 44587 -2250
rect 26779 -2314 44587 -2268
rect 47973 -1786 68149 -1760
rect 47973 -1830 67596 -1786
rect 47973 -2172 48050 -1830
rect 48308 -2172 67596 -1830
rect 47973 -2272 67596 -2172
rect 68018 -2272 68149 -1786
rect 47973 -2314 68149 -2272
rect 71635 -1830 91015 -1760
rect 71635 -2146 71670 -1830
rect 71936 -1876 91015 -1830
rect 71936 -2146 90546 -1876
rect 71635 -2244 90546 -2146
rect 90922 -2244 91015 -1876
rect 71635 -2314 91015 -2244
rect 94575 -1804 117458 -1760
rect 94575 -2230 94660 -1804
rect 94952 -2230 117458 -1804
rect 94575 -2314 117458 -2230
rect 11892 -2320 11964 -2314
rect 17014 -2315 17084 -2314
rect 20212 -2316 20274 -2314
rect 26990 -2316 27382 -2314
rect 27954 -2322 28026 -2314
rect 58636 -2318 58708 -2314
rect 67212 -2315 67278 -2314
rect 19004 -2722 20346 -2622
rect 19004 -3184 19172 -2722
rect 20150 -3184 20346 -2722
rect 19004 -3278 20346 -3184
rect 42944 -2686 44082 -2606
rect 42944 -3226 43016 -2686
rect 43986 -3226 44082 -2686
rect 42944 -3268 44082 -3226
rect 65758 -2732 67080 -2618
rect 65758 -3166 65848 -2732
rect 66898 -3166 67080 -2732
rect 65758 -3258 67080 -3166
rect 89696 -2722 91328 -2626
rect 89696 -3208 89834 -2722
rect 91108 -3208 91328 -2722
rect 89696 -3304 91328 -3208
rect 26394 -3990 27668 -3868
rect 26394 -4446 26522 -3990
rect 27568 -4446 27668 -3990
rect 26394 -4526 27668 -4446
rect 50940 -3928 51898 -3874
rect 50940 -4472 51026 -3928
rect 51844 -4472 51898 -3928
rect 50940 -4526 51898 -4472
rect 73315 -4010 75340 -3886
rect 73315 -4448 73494 -4010
rect 75202 -4448 75340 -4010
rect 73315 -4529 75340 -4448
rect 97388 -4008 99380 -3886
rect 97388 -4410 97540 -4008
rect 99214 -4410 99380 -4008
rect 97388 -4522 99380 -4410
<< via3 >>
rect 19172 -3184 20150 -2722
rect 43016 -3226 43986 -2686
rect 65848 -3166 66898 -2732
rect 89834 -3208 91108 -2722
rect 26522 -4446 27568 -3990
rect 51026 -4472 51844 -3928
rect 73494 -4448 75202 -4010
rect 97540 -4410 99214 -4008
<< metal4 >>
rect 878 -2617 1536 4073
rect 39957 -2617 40655 2817
rect 42944 -2617 44082 -2606
rect 53908 -2617 54559 3171
rect 85999 -2617 86697 2807
rect 102481 -2617 103139 2975
rect 878 -2686 103139 -2617
rect 878 -2722 43016 -2686
rect 878 -3184 19172 -2722
rect 20150 -3184 43016 -2722
rect 878 -3226 43016 -3184
rect 43986 -2722 103139 -2686
rect 43986 -2732 89834 -2722
rect 43986 -3166 65848 -2732
rect 66898 -3166 89834 -2732
rect 43986 -3208 89834 -3166
rect 91108 -3208 103139 -2722
rect 43986 -3226 103139 -3208
rect 878 -3275 103139 -3226
rect 19004 -3278 20346 -3275
rect 85999 -3399 86697 -3275
rect 26394 -3990 27668 -3868
rect 26394 -4446 26522 -3990
rect 27568 -4446 27668 -3990
rect 26394 -4526 27668 -4446
rect 50940 -3928 51898 -3874
rect 50940 -4472 51026 -3928
rect 51844 -4472 51898 -3928
rect 50940 -4526 51898 -4472
rect 73315 -4010 75340 -3886
rect 73315 -4448 73494 -4010
rect 75202 -4448 75340 -4010
rect 73315 -4529 75340 -4448
rect 97388 -4008 99380 -3886
rect 97388 -4410 97540 -4008
rect 99214 -4410 99380 -4008
rect 97388 -4522 99380 -4410
<< via4 >>
rect 26522 -4446 27568 -3990
rect 51026 -4472 51844 -3928
rect 73494 -4448 75202 -4010
rect 97540 -4410 99214 -4008
<< metal5 >>
rect 284 -3871 942 8622
rect 15989 -3871 16647 3185
rect 31459 -3871 32117 2977
rect 62187 -3871 62845 3079
rect 77709 -3871 78367 2967
rect 116571 -3871 117161 4771
rect 284 -3928 117161 -3871
rect 284 -3990 51026 -3928
rect 284 -4446 26522 -3990
rect 27568 -4446 51026 -3990
rect 284 -4472 51026 -4446
rect 51844 -4008 117161 -3928
rect 51844 -4010 97540 -4008
rect 51844 -4448 73494 -4010
rect 75202 -4410 97540 -4010
rect 99214 -4410 117161 -4008
rect 75202 -4448 117161 -4410
rect 51844 -4472 117161 -4448
rect 284 -4529 117161 -4472
rect 116571 -4599 117161 -4529
use buffer_digital  buffer_digital_0 ~/Desktop/charge_pumps2/layout_files
timestamp 1698753667
transform 1 0 20636 0 1 -2364
box -274 0 415 576
use buffer_digital  buffer_digital_1
timestamp 1698753667
transform 1 0 26404 0 1 -2348
box -274 0 415 576
use buffer_digital  buffer_digital_2
timestamp 1698753667
transform 1 0 44680 0 1 -2276
box -274 0 415 576
use buffer_digital  buffer_digital_3
timestamp 1698753667
transform 1 0 47556 0 1 -2286
box -274 0 415 576
use buffer_digital  buffer_digital_4
timestamp 1698753667
transform 1 0 68218 0 1 -2230
box -274 0 415 576
use buffer_digital  buffer_digital_5
timestamp 1698753667
transform 1 0 71218 0 1 -2216
box -274 0 415 576
use buffer_digital  buffer_digital_6
timestamp 1698753667
transform 1 0 91076 0 1 -2312
box -274 0 415 576
use buffer_digital  buffer_digital_7
timestamp 1698753667
transform 1 0 94166 0 1 -2290
box -274 0 415 576
use charge_pump  charge_pump_0
timestamp 1698757234
transform 1 0 -480 0 1 7870
box 498 -7862 23756 19014
use charge_pump  charge_pump_1
timestamp 1698757234
transform 1 0 46226 0 1 7872
box 498 -7862 23756 19014
use charge_pump  charge_pump_2
timestamp 1698757234
transform 1 0 93528 0 1 7864
box 498 -7862 23756 19014
use charge_pump_reverse  charge_pump_reverse_0
timestamp 1698753667
transform 1 0 22894 0 -1 24894
box 498 -3206 23756 25968
use charge_pump_reverse  charge_pump_reverse_1
timestamp 1698753667
transform 1 0 69556 0 -1 24884
box 498 -3206 23756 25968
<< end >>
