magic
tech sky130A
magscale 1 2
timestamp 1699075837
<< nwell >>
rect 3128 308 6366 888
rect 7840 300 8660 626
rect 10938 306 13150 890
rect 22878 192 25166 764
<< nsubdiff >>
rect 8012 524 8190 548
rect 8012 370 8038 524
rect 8154 370 8190 524
rect 8012 352 8190 370
<< nsubdiffcont >>
rect 8038 370 8154 524
<< locali >>
rect 8012 524 8190 548
rect 8012 370 8038 524
rect 8154 370 8190 524
rect 8012 352 8190 370
<< viali >>
rect 8038 370 8154 524
<< metal1 >>
rect 23559 26724 23927 27196
rect 23659 26688 23927 26724
rect 832 7360 1272 9514
rect 832 6628 936 7360
rect 1120 6628 1272 7360
rect 832 1002 1272 6628
rect 1578 7420 2006 7432
rect 1578 7348 2020 7420
rect 1578 6432 1674 7348
rect 1938 6432 2020 7348
rect 1578 6380 2020 6432
rect 1578 1052 2006 6380
rect 24656 1052 25052 7154
rect 832 540 1290 1002
rect 1578 994 25052 1052
rect 1578 808 7532 994
rect 8980 808 25052 994
rect 1578 650 25052 808
rect 1600 644 24906 650
rect 7450 600 9094 644
rect 8036 548 8156 600
rect 846 -12 1290 540
rect 8012 524 8190 548
rect 1930 -12 6418 428
rect 8012 370 8038 524
rect 8154 370 8190 524
rect 8012 352 8190 370
rect 9154 386 9514 422
rect 9154 252 9188 386
rect 7768 199 8520 232
rect 9016 219 9188 252
rect 7460 -10 7494 86
rect 7678 -10 7712 86
rect 8706 36 8740 102
rect 8924 36 8958 102
rect 9154 88 9188 219
rect 9462 88 9514 386
rect 9154 56 9514 88
rect 8706 12 8958 36
rect 8652 -10 9018 12
rect 7456 -12 9018 -10
rect 9854 -12 13168 440
rect 14776 -12 21690 394
rect 21932 -12 25160 302
rect 25362 -12 25808 7960
rect 846 -56 25808 -12
rect 846 -262 7522 -56
rect 8864 -262 25808 -56
rect 846 -404 25808 -262
rect 846 -408 25758 -404
rect 932 -446 25758 -408
<< via1 >>
rect 936 6628 1120 7360
rect 1674 6432 1938 7348
rect 7532 808 8980 994
rect 9188 88 9462 386
rect 7522 -262 8864 -56
<< metal2 >>
rect 870 7360 1190 7482
rect 870 6628 936 7360
rect 1120 6628 1190 7360
rect 870 6562 1190 6628
rect 1578 7348 2020 7420
rect 1578 6432 1674 7348
rect 1938 6432 2020 7348
rect 1578 6380 2020 6432
rect 7458 1046 7818 1048
rect 7458 994 9078 1046
rect 7458 808 7532 994
rect 8980 808 9078 994
rect 7458 756 9078 808
rect 7458 748 7818 756
rect 6586 402 7258 426
rect 6586 78 6648 402
rect 7052 317 7258 402
rect 9154 386 9514 422
rect 7052 111 7391 317
rect 7052 78 7258 111
rect 6586 52 7258 78
rect 9154 88 9188 386
rect 9462 88 9514 386
rect 9154 56 9514 88
rect 7456 -56 8966 -10
rect 7456 -262 7522 -56
rect 8864 -262 8966 -56
rect 7456 -302 8966 -262
<< via2 >>
rect 936 6628 1120 7360
rect 1674 6432 1938 7348
rect 7532 808 8980 994
rect 6648 78 7052 402
rect 9188 88 9462 386
rect 7522 -262 8864 -56
<< metal3 >>
rect 870 7360 1190 7482
rect 870 6628 936 7360
rect 1120 6628 1190 7360
rect 870 6562 1190 6628
rect 1578 7348 2020 7420
rect 1578 6432 1674 7348
rect 1938 6432 2020 7348
rect 1578 6380 2020 6432
rect 13346 1140 13418 1642
rect 7458 1046 7818 1048
rect 7458 994 9078 1046
rect 7458 808 7532 994
rect 8980 808 9078 994
rect 7458 756 9078 808
rect 7458 748 7818 756
rect 6586 424 7258 426
rect 13297 424 13431 1140
rect 1805 402 7258 424
rect 1805 78 6648 402
rect 7052 78 7258 402
rect 1805 52 7258 78
rect 9144 386 25666 424
rect 9144 88 9188 386
rect 9462 332 25666 386
rect 9462 88 25447 332
rect 1805 46 6916 52
rect 9144 46 25447 88
rect 7456 -56 8966 -10
rect 7456 -262 7522 -56
rect 8864 -262 8966 -56
rect 7456 -302 8966 -262
<< via3 >>
rect 936 6628 1120 7360
rect 1674 6432 1938 7348
rect 7532 808 8980 994
rect 7522 -262 8864 -56
<< metal4 >>
rect 870 7360 1190 7482
rect 870 6628 936 7360
rect 1182 6628 1190 7360
rect 870 6562 1190 6628
rect 1488 7348 2056 12518
rect 1488 6432 1674 7348
rect 1938 6432 2056 7348
rect 1488 1136 2056 6432
rect 24592 1136 25160 7494
rect 1488 994 25160 1136
rect 1488 808 7532 994
rect 8980 808 25160 994
rect 1488 578 25160 808
rect 1488 568 24670 578
rect 7456 -28 8966 -10
rect 7456 -276 7518 -28
rect 8874 -276 8966 -28
rect 7456 -302 8966 -276
<< via4 >>
rect 936 6628 1120 7360
rect 1120 6628 1182 7360
rect 7518 -56 8874 -28
rect 7518 -262 7522 -56
rect 7522 -262 8864 -56
rect 8864 -262 8874 -56
rect 7518 -276 8874 -262
<< metal5 >>
rect 789 7360 1393 10802
rect 789 6628 936 7360
rect 1182 6628 1393 7360
rect 789 46 1393 6628
rect 25314 46 25904 10915
rect 789 -28 25904 46
rect 789 -276 7518 -28
rect 8874 -276 25904 -28
rect 789 -507 25904 -276
rect 789 -558 25892 -507
use buffer_digital  buffer_digital_0
timestamp 1699074083
transform 1 0 8708 0 1 68
box -274 -74 412 576
use buffer_digital  buffer_digital_1
timestamp 1699074083
transform 1 0 7462 0 1 52
box -274 -74 412 576
use charge_pump1_reverse  charge_pump1_reverse_0
timestamp 1699075837
transform 1 0 821 0 -1 27108
box -313 -2944 25321 25896
use nmos_decap_10  nmos_decap_10_0
timestamp 1698837560
transform 0 1 1262 -1 0 2080
box -10 -42 1060 416
use nmos_decap_10  nmos_decap_10_1
timestamp 1698837560
transform 0 1 1262 -1 0 3040
box -10 -42 1060 416
use nmos_decap_10  nmos_decap_10_2
timestamp 1698837560
transform 0 1 1262 -1 0 4000
box -10 -42 1060 416
use nmos_decap_10  nmos_decap_10_3
timestamp 1698837560
transform 0 1 1262 -1 0 4960
box -10 -42 1060 416
use nmos_decap_10  nmos_decap_10_4
timestamp 1698837560
transform 0 1 1262 -1 0 5920
box -10 -42 1060 416
use nmos_decap_10  nmos_decap_10_5
timestamp 1698837560
transform 1 0 13860 0 1 352
box -10 -42 1060 416
use nmos_decap_10  nmos_decap_10_6
timestamp 1698837560
transform 1 0 14820 0 1 352
box -10 -42 1060 416
use nmos_decap_10  nmos_decap_10_7
timestamp 1698837560
transform 1 0 15780 0 1 352
box -10 -42 1060 416
use nmos_decap_10  nmos_decap_10_8
timestamp 1698837560
transform 1 0 16740 0 1 352
box -10 -42 1060 416
use nmos_decap_10  nmos_decap_10_9
timestamp 1698837560
transform 1 0 17700 0 1 352
box -10 -42 1060 416
use nmos_decap_10  nmos_decap_10_10
timestamp 1698837560
transform 1 0 18660 0 1 352
box -10 -42 1060 416
use nmos_decap_10  nmos_decap_10_11
timestamp 1698837560
transform 1 0 19620 0 1 352
box -10 -42 1060 416
use nmos_decap_10  nmos_decap_10_12
timestamp 1698837560
transform 1 0 20580 0 1 352
box -10 -42 1060 416
use pmos_decap_10  pmos_decap_10_0
timestamp 1698841269
transform 0 1 25002 -1 0 2222
box 0 -108 1098 464
use pmos_decap_10  pmos_decap_10_1
timestamp 1698841269
transform 0 1 25006 -1 0 3572
box 0 -108 1098 464
use pmos_decap_10  pmos_decap_10_2
timestamp 1698841269
transform 0 1 25006 -1 0 4920
box 0 -108 1098 464
use pmos_decap_10  pmos_decap_10_3
timestamp 1698841269
transform 0 1 25022 -1 0 6270
box 0 -108 1098 464
use pmos_decap_10  pmos_decap_10_4
timestamp 1698841269
transform 0 1 25044 -1 0 7660
box 0 -108 1098 464
use pmos_decap_10  pmos_decap_10_5
timestamp 1698841269
transform 1 0 2056 0 -1 770
box 0 -108 1098 464
use pmos_decap_10  pmos_decap_10_6
timestamp 1698841269
transform 1 0 3128 0 -1 772
box 0 -108 1098 464
use pmos_decap_10  pmos_decap_10_7
timestamp 1698841269
transform 1 0 4200 0 -1 772
box 0 -108 1098 464
use pmos_decap_10  pmos_decap_10_8
timestamp 1698841269
transform 1 0 5272 0 -1 778
box 0 -108 1098 464
use pmos_decap_10  pmos_decap_10_9
timestamp 1698841269
transform 1 0 9896 0 -1 768
box 0 -108 1098 464
use pmos_decap_10  pmos_decap_10_10
timestamp 1698841269
transform 1 0 10968 0 -1 774
box 0 -108 1098 464
use pmos_decap_10  pmos_decap_10_11
timestamp 1698841269
transform 1 0 12042 0 -1 774
box 0 -108 1098 464
use pmos_decap_10  pmos_decap_10_12
timestamp 1698841269
transform 1 0 21932 0 -1 652
box 0 -108 1098 464
use pmos_decap_10  pmos_decap_10_13
timestamp 1698841269
transform 1 0 23004 0 -1 662
box 0 -108 1098 464
use pmos_decap_10  pmos_decap_10_14
timestamp 1698841269
transform 1 0 24076 0 -1 666
box 0 -108 1098 464
<< end >>
