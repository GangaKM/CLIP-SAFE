magic
tech sky130A
magscale 1 2
timestamp 1698902493
<< nwell >>
rect 0 242 992 502
rect 0 0 930 242
rect -32 -498 930 -288
rect -32 -858 978 -498
<< nsubdiff >>
rect 186 434 282 460
rect 186 398 216 434
rect 254 398 282 434
rect 186 372 282 398
rect 846 -706 942 -680
rect 846 -742 876 -706
rect 914 -742 942 -706
rect 846 -768 942 -742
<< nsubdiffcont >>
rect 216 398 254 434
rect 876 -742 914 -706
<< locali >>
rect 186 442 282 460
rect 186 392 202 442
rect 266 392 282 442
rect 186 372 282 392
rect 846 -698 942 -680
rect 846 -748 862 -698
rect 926 -748 942 -698
rect 846 -768 942 -748
<< viali >>
rect -54 524 1000 586
rect 202 434 266 442
rect 202 398 216 434
rect 216 398 254 434
rect 254 398 266 434
rect 202 392 266 398
rect 862 -706 926 -698
rect 862 -742 876 -706
rect 876 -742 914 -706
rect 914 -742 926 -706
rect 862 -748 926 -742
rect -34 -1022 974 -908
<< metal1 >>
rect -66 586 1020 616
rect -66 524 -54 586
rect 1000 524 1020 586
rect -66 498 1020 524
rect 50 436 84 498
rect 246 448 276 460
rect 190 442 278 448
rect 190 436 202 442
rect 50 392 202 436
rect 266 392 278 442
rect 50 388 278 392
rect 50 110 84 388
rect 190 386 278 388
rect 880 242 952 292
rect 880 130 938 242
rect 864 16 938 130
rect 20 -530 70 -364
rect 20 -600 92 -530
rect 884 -548 938 16
rect 20 -646 108 -600
rect 20 -788 92 -646
rect 906 -692 936 -548
rect 850 -698 938 -692
rect 850 -748 862 -698
rect 926 -748 938 -698
rect 850 -754 938 -748
rect -38 -902 984 -788
rect -46 -908 986 -902
rect -46 -1022 -34 -908
rect 974 -1022 986 -908
rect -46 -1028 986 -1022
rect -38 -1120 984 -1028
<< via1 >>
rect -54 524 1000 586
rect -34 -1022 974 -908
<< metal2 >>
rect -66 586 1020 616
rect -66 524 -54 586
rect 1000 524 1020 586
rect -66 498 1020 524
rect -38 -908 984 -788
rect -38 -1022 -34 -908
rect 974 -1022 984 -908
rect -38 -1120 984 -1022
<< via2 >>
rect -54 524 1000 586
rect -34 -1022 974 -908
<< metal3 >>
rect -64 524 -54 594
rect 1006 524 1016 594
rect -64 519 1010 524
rect -38 -820 984 -788
rect -48 -836 -38 -820
rect -52 -1050 -42 -836
rect -48 -1088 -38 -1050
rect 984 -1088 994 -820
rect -38 -1120 984 -1088
<< via3 >>
rect -54 586 1006 594
rect -54 524 1000 586
rect 1000 524 1006 586
rect -38 -836 984 -820
rect -42 -908 984 -836
rect -42 -1022 -34 -908
rect -34 -1022 974 -908
rect 974 -1022 984 -908
rect -42 -1050 984 -1022
rect -38 -1088 984 -1050
<< metal4 >>
rect -62 616 1022 620
rect -66 594 1022 616
rect -66 524 -54 594
rect 1006 524 1022 594
rect -66 500 1022 524
rect -66 498 1020 500
rect -38 -819 984 -788
rect -39 -820 985 -819
rect -39 -835 -38 -820
rect -43 -836 -38 -835
rect -43 -1050 -42 -836
rect -43 -1051 -38 -1050
rect -39 -1088 -38 -1051
rect 984 -1088 985 -820
rect -39 -1089 985 -1088
rect -38 -1120 984 -1089
<< via4 >>
rect -38 -1088 984 -820
<< metal5 >>
rect -62 -820 1008 -786
rect -62 -1088 -38 -820
rect 984 -1088 1008 -820
rect -62 -1112 1008 -1088
rect -38 -1120 984 -1112
use sky130_fd_pr__pfet_01v8_lvt_46RJ2R  sky130_fd_pr__pfet_01v8_lvt_46RJ2R_0
timestamp 1698771642
transform 1 0 494 0 1 164
box -494 -164 494 198
use sky130_fd_pr__pfet_01v8_lvt_46RJ2R  sky130_fd_pr__pfet_01v8_lvt_46RJ2R_1
timestamp 1698771642
transform 1 0 480 0 1 -490
box -494 -164 494 198
<< labels >>
rlabel metal4 544 612 544 612 1 Vdd
port 1 n
rlabel metal5 470 -1100 470 -1100 1 gnd
port 2 n
rlabel metal1 900 -144 900 -144 1 vout
<< end >>
