magic
tech sky130A
magscale 1 2
timestamp 1698152391
<< nwell >>
rect 1358 2036 1492 2084
rect 1426 2032 1492 2036
rect 1468 1640 1492 2032
<< poly >>
rect 206 2074 236 2078
rect -1140 2042 1390 2074
rect -1138 1994 -1108 2042
rect -946 1994 -916 2042
rect -754 1994 -724 2042
rect -562 1996 -532 2042
rect -370 1994 -340 2042
rect -178 1998 -148 2042
rect 14 1996 44 2042
rect 206 2002 236 2042
rect 398 1994 428 2042
rect 590 1998 620 2042
rect 782 1998 812 2042
rect 974 1998 1004 2042
rect 1166 1998 1196 2042
rect 1358 1996 1388 2042
rect -1138 1692 -1108 1725
rect -1042 1692 -1012 1736
rect -850 1692 -820 1736
rect -658 1692 -628 1736
rect -466 1692 -436 1736
rect -274 1692 -244 1738
rect -82 1692 -52 1736
rect 110 1692 140 1736
rect 302 1692 332 1738
rect 494 1692 524 1736
rect 686 1692 716 1738
rect 878 1692 908 1736
rect 1070 1692 1100 1736
rect 1262 1692 1292 1736
rect 1358 1692 1388 1695
rect -1158 1658 1391 1692
rect -1138 1555 -1108 1658
rect 1357 1640 1391 1658
rect 1358 1578 1388 1640
rect -562 1555 -532 1556
rect 974 1555 1004 1556
rect 1166 1555 1196 1556
rect 1357 1555 1391 1578
rect -1139 1521 1391 1555
rect -1138 1482 -1108 1521
rect -946 1484 -916 1521
rect -754 1486 -724 1521
rect -562 1488 -532 1521
rect -370 1486 -340 1521
rect -178 1486 -148 1521
rect 14 1486 44 1521
rect 206 1486 236 1521
rect 398 1486 428 1521
rect 590 1486 620 1521
rect 782 1484 812 1521
rect 974 1488 1004 1521
rect 1166 1488 1196 1521
rect 1358 1488 1388 1521
rect -1042 1360 -1012 1398
rect -850 1360 -820 1398
rect -658 1360 -628 1398
rect -466 1360 -436 1408
rect -274 1360 -244 1398
rect -82 1360 -52 1396
rect 110 1360 140 1394
rect 302 1360 332 1394
rect 494 1360 524 1394
rect 686 1360 716 1394
rect 878 1360 908 1398
rect 1070 1360 1100 1394
rect 1262 1360 1292 1396
rect -1157 1326 1406 1360
<< locali >>
rect -1061 2072 1390 2074
rect -1140 2040 1390 2072
rect -1140 2038 -1044 2040
rect 1228 2038 1310 2040
rect -1156 1658 1390 1694
rect 1354 1556 1390 1658
rect -1138 1520 1390 1556
rect -1156 1324 1406 1360
<< metal1 >>
rect -1188 2110 1347 2140
rect -1188 1912 -1154 2110
rect -1104 1980 -1046 1992
rect -1048 1752 -1046 1980
rect -996 1908 -962 2110
rect -914 1980 -856 1992
rect -1104 1740 -1046 1752
rect -914 1752 -912 1980
rect -804 1918 -770 2110
rect -718 1980 -660 1992
rect -914 1740 -856 1752
rect -662 1752 -660 1980
rect -612 1916 -578 2110
rect -526 1980 -468 1992
rect -718 1740 -660 1752
rect -470 1752 -468 1980
rect -420 1920 -386 2110
rect -336 1980 -278 1992
rect -526 1740 -468 1752
rect -280 1752 -278 1980
rect -228 1914 -194 2110
rect -144 1980 -86 1992
rect -336 1740 -278 1752
rect -144 1752 -142 1980
rect -36 1912 -2 2110
rect 48 1980 106 1992
rect -144 1740 -86 1752
rect 48 1752 50 1980
rect 156 1912 190 2110
rect 240 1980 298 1992
rect 48 1740 106 1752
rect 296 1752 298 1980
rect 348 1908 382 2110
rect 432 1980 490 1994
rect 240 1740 298 1752
rect 488 1752 490 1980
rect 540 1904 574 2110
rect 626 1980 684 1994
rect 432 1742 490 1752
rect 682 1752 684 1980
rect 732 1918 766 2110
rect 816 1980 874 1992
rect 626 1742 684 1752
rect 816 1752 818 1980
rect 924 1870 958 2110
rect 1008 1980 1066 1992
rect 816 1740 874 1752
rect 1064 1752 1066 1980
rect 1116 1874 1150 2110
rect 1200 1980 1258 1992
rect 1008 1740 1066 1752
rect 1256 1752 1258 1980
rect 1317 1753 1347 2110
rect 1392 1980 1452 1992
rect 1200 1740 1258 1752
rect 1392 1752 1394 1980
rect 1450 1752 1452 1980
rect 1392 1742 1452 1752
rect 1404 1738 1444 1742
rect 1408 1612 1444 1738
rect 1306 1576 1512 1612
rect -1102 1470 -1044 1484
rect -1188 1398 -1154 1438
rect -1046 1410 -1044 1470
rect -910 1470 -852 1484
rect -1102 1398 -1044 1410
rect -996 1398 -962 1432
rect -854 1410 -852 1470
rect -720 1470 -662 1484
rect -910 1398 -852 1410
rect -804 1398 -770 1428
rect -664 1410 -662 1470
rect -528 1470 -470 1484
rect -720 1398 -662 1410
rect -612 1398 -578 1434
rect -472 1410 -470 1470
rect -338 1470 -280 1484
rect -528 1398 -470 1410
rect -420 1398 -386 1432
rect -338 1410 -336 1470
rect -144 1470 -86 1484
rect -338 1398 -280 1410
rect -228 1398 -194 1434
rect -88 1410 -86 1470
rect 48 1470 106 1484
rect -144 1398 -86 1410
rect -36 1398 -2 1432
rect 104 1410 106 1470
rect 242 1470 300 1484
rect 48 1398 106 1410
rect 156 1398 190 1430
rect 298 1410 300 1470
rect 434 1470 492 1484
rect 242 1398 300 1410
rect 348 1398 382 1436
rect 490 1410 492 1470
rect 624 1470 682 1484
rect 434 1398 492 1410
rect 540 1398 574 1434
rect 680 1410 682 1470
rect 818 1470 876 1484
rect 624 1398 682 1410
rect 732 1398 766 1432
rect 874 1410 876 1470
rect 1008 1470 1066 1484
rect 818 1398 876 1410
rect 924 1398 958 1434
rect 1064 1410 1066 1470
rect 1200 1470 1258 1484
rect 1008 1398 1066 1410
rect 1116 1398 1150 1434
rect 1256 1410 1258 1470
rect 1306 1430 1342 1576
rect 1404 1484 1438 1488
rect 1392 1470 1450 1484
rect 1200 1398 1258 1410
rect 1309 1398 1343 1423
rect 1448 1410 1450 1470
rect 1392 1398 1450 1410
<< via1 >>
rect -1104 1752 -1048 1980
rect -912 1752 -856 1980
rect -718 1752 -662 1980
rect -526 1752 -470 1980
rect -336 1752 -280 1980
rect -142 1752 -86 1980
rect 50 1752 106 1980
rect 240 1752 296 1980
rect 432 1752 488 1980
rect 626 1752 682 1980
rect 818 1752 874 1980
rect 1008 1752 1064 1980
rect 1200 1752 1256 1980
rect 1394 1752 1450 1980
rect -1102 1410 -1046 1470
rect -910 1410 -854 1470
rect -720 1410 -664 1470
rect -528 1410 -472 1470
rect -336 1410 -280 1470
rect -144 1410 -88 1470
rect 48 1410 104 1470
rect 242 1410 298 1470
rect 434 1410 490 1470
rect 624 1410 680 1470
rect 818 1410 874 1470
rect 1008 1410 1064 1470
rect 1200 1410 1256 1470
rect 1392 1410 1448 1470
<< metal2 >>
rect -1144 1980 1450 1992
rect -1144 1752 -1104 1980
rect -1048 1752 -912 1980
rect -856 1752 -718 1980
rect -662 1752 -526 1980
rect -470 1752 -336 1980
rect -280 1752 -142 1980
rect -86 1752 50 1980
rect 106 1752 240 1980
rect 296 1752 432 1980
rect 488 1752 626 1980
rect 682 1752 818 1980
rect 874 1752 1008 1980
rect 1064 1752 1200 1980
rect 1256 1752 1394 1980
rect -1144 1740 1450 1752
rect -1138 1470 1450 1484
rect -1138 1410 -1102 1470
rect -1046 1410 -910 1470
rect -854 1410 -720 1470
rect -664 1410 -528 1470
rect -472 1410 -336 1470
rect -280 1410 -144 1470
rect -88 1410 48 1470
rect 104 1410 242 1470
rect 298 1410 434 1470
rect 490 1410 624 1470
rect 680 1410 818 1470
rect 874 1410 1008 1470
rect 1064 1410 1200 1470
rect 1256 1410 1392 1470
rect 1448 1410 1450 1470
rect -1138 1398 1450 1410
use sky130_fd_pr__nfet_01v8_NJGLN5  sky130_fd_pr__nfet_01v8_NJGLN5_1 ~/Desktop/charge_pumps2/layout_files
timestamp 1698060067
transform 1 0 125 0 1 1440
box -1325 -130 1325 130
use sky130_fd_pr__pfet_01v8_VR4B8J  sky130_fd_pr__pfet_01v8_VR4B8J_1 ~/Desktop/charge_pumps2/layout_files
timestamp 1698060067
transform 1 0 125 0 1 1858
box -1361 -226 1361 226
<< end >>
