magic
tech sky130A
magscale 1 2
timestamp 1699075837
<< error_p >>
rect 57471 25408 57479 25410
rect 57499 25408 57507 25410
rect 20045 25402 20053 25404
rect 20073 25402 20081 25404
rect 71869 25398 71877 25400
rect 71897 25398 71905 25400
rect 20037 23310 20045 23312
rect 20065 23310 20073 23312
rect 71861 23306 71869 23308
rect 71889 23306 71897 23308
rect 57441 23302 57449 23304
rect 57469 23302 57477 23304
rect 71837 21212 71845 21214
rect 71865 21212 71873 21214
rect 57445 21208 57453 21210
rect 57473 21208 57481 21210
<< metal2 >>
rect 51697 27705 51863 28213
rect 103241 28104 103828 28188
rect 51697 27539 51990 27705
rect 103744 27538 103828 28104
rect 23904 26322 28100 26408
rect 50126 26372 53544 26456
rect 75752 26356 79622 26450
rect 101678 26346 105512 26408
rect 23920 24230 28116 24316
rect 50134 24278 53552 24362
rect 75748 24266 79618 24360
rect 101674 24264 105468 24304
rect 23886 22142 28082 22228
rect 50166 22184 53584 22268
rect 75690 22160 79600 22224
rect 101700 22158 105410 22208
rect 23938 20058 28100 20170
rect 50214 20098 53552 20174
rect 75774 20064 79722 20124
rect 101758 20072 105468 20122
rect 23894 17968 28056 18080
rect 50246 18002 53584 18078
rect 75730 17974 79678 18034
rect 101802 17986 105518 18020
rect 23816 15828 28084 15936
rect 50204 15908 53580 16012
rect 75662 15874 79610 15934
rect 101736 15882 105506 15928
rect 23820 13764 28086 13834
rect 50248 13826 53586 13882
rect 75642 13790 79590 13850
rect 101772 13800 105538 13834
rect 23820 11670 28114 11742
rect 50242 11714 53626 11778
rect 75664 11678 79648 11756
rect 101790 11700 105556 11734
rect 26256 9994 26340 10598
rect 25393 9910 26340 9994
rect 77818 9990 77902 10564
rect 77217 9906 77902 9990
<< metal3 >>
rect 8678 604 32823 982
rect 8678 572 28091 604
rect 35015 600 58418 978
rect 75934 852 84560 978
rect 8678 502 9024 572
rect 10388 502 28091 572
rect 50352 502 58418 600
rect 60505 474 84560 852
rect 102127 474 110361 852
<< metal4 >>
rect -578 27464 -10 27474
rect -578 26888 12394 27464
rect 116994 26890 129854 27466
rect -578 25350 -10 26888
rect 129236 25352 129804 26890
rect -578 24796 12159 25350
rect 115389 24798 129804 25352
rect -578 23258 -10 24796
rect 129236 23260 129804 24798
rect -578 22704 12159 23258
rect 117307 22706 129804 23260
rect -578 21158 -10 22704
rect 129236 21160 129804 22706
rect -578 20604 12273 21158
rect 117219 20606 129804 21160
rect -578 19088 -10 20604
rect 129236 19090 129804 20606
rect -578 18544 12222 19088
rect 117224 18546 129804 19090
rect -578 16978 -10 18544
rect 129236 16980 129804 18546
rect -578 16434 12312 16978
rect 117246 16436 129804 16980
rect -578 14894 -10 16434
rect 129236 14910 129804 16436
rect -578 14364 12215 14894
rect 117136 14366 129804 14910
rect -578 12776 -10 14364
rect 129236 12778 129804 14366
rect -578 12232 12222 12776
rect 117202 12234 129804 12778
rect -578 5506 -10 12232
rect -622 4938 7364 5506
rect -578 1694 -10 4938
rect -578 1126 4214 1694
rect 24084 1136 27838 1704
rect 50412 1142 53584 1690
rect 50412 1122 52056 1142
rect 52772 1122 53584 1142
rect 75908 1132 79384 1700
rect 129236 1696 129804 12234
rect 101988 1154 105372 1696
rect 101988 1128 103924 1154
rect 104724 1128 105372 1154
rect 122968 1128 129804 1696
<< metal5 >>
rect -1312 28542 2086 29146
rect -1312 25992 -708 28542
rect -1312 25416 12234 25992
rect 117996 25909 130440 25994
rect 117996 25418 130459 25909
rect -1312 23864 -708 25416
rect 304 25106 356 25416
rect 129869 23866 130459 25418
rect -1312 23310 12201 23864
rect 119227 23312 130459 23866
rect -1312 21774 -708 23310
rect 129869 21776 130459 23312
rect -1331 21220 12179 21774
rect 119193 21222 130459 21776
rect -1312 19674 -708 21220
rect 129869 19676 130459 21222
rect -1312 19130 12152 19674
rect 119242 19132 130524 19676
rect -1312 17604 -708 19130
rect 129869 17606 130459 19132
rect -1312 17060 12218 17604
rect 118732 17062 130459 17606
rect -1312 15514 -708 17060
rect 129869 15516 130459 17062
rect -1312 14970 12152 15514
rect 118800 14972 130459 15516
rect -1312 13434 -708 14970
rect 129869 13436 130459 14972
rect -1312 12890 12218 13434
rect 118944 12892 130459 13436
rect -1312 604 -708 12890
rect 129869 5869 130459 12892
rect 125221 5279 130459 5869
rect -1312 0 6420 604
rect 24646 0 27410 604
rect 51124 -4 52709 600
rect 76558 -4 78736 600
rect 102674 2 104712 606
use cp1_buffer1  cp1_buffer1_0
timestamp 1699075837
transform 1 0 -508 0 1 558
box 508 -558 26142 29136
use cp1_buffer1  cp1_buffer1_1
timestamp 1699075837
transform 1 0 51316 0 1 554
box 508 -558 26142 29136
use cp1_buffer1  cp1_buffer1_2
timestamp 1699075837
transform 1 0 103260 0 1 560
box 508 -558 26142 29136
use cp1_buffer1_reverse  cp1_buffer1_reverse_0
timestamp 1699075837
transform 1 0 25806 0 1 456
box 508 -558 26142 30052
use cp1_buffer1_reverse  cp1_buffer1_reverse_1
timestamp 1699075837
transform 1 0 77340 0 1 428
box 508 -558 26142 30052
<< end >>
