magic
tech sky130A
magscale 1 2
timestamp 1697701953
<< nwell >>
rect -257 188 353 226
rect -353 -188 353 188
rect -353 -226 257 -188
<< pmos >>
rect -255 -126 -225 126
rect -159 -126 -129 126
rect -63 -126 -33 126
rect 33 -126 63 126
rect 129 -126 159 126
rect 225 -126 255 126
<< pdiff >>
rect -317 114 -255 126
rect -317 -114 -305 114
rect -271 -114 -255 114
rect -317 -126 -255 -114
rect -225 114 -159 126
rect -225 -114 -209 114
rect -175 -114 -159 114
rect -225 -126 -159 -114
rect -129 114 -63 126
rect -129 -114 -113 114
rect -79 -114 -63 114
rect -129 -126 -63 -114
rect -33 114 33 126
rect -33 -114 -17 114
rect 17 -114 33 114
rect -33 -126 33 -114
rect 63 114 129 126
rect 63 -114 79 114
rect 113 -114 129 114
rect 63 -126 129 -114
rect 159 114 225 126
rect 159 -114 175 114
rect 209 -114 225 114
rect 159 -126 225 -114
rect 255 114 317 126
rect 255 -114 271 114
rect 305 -114 317 114
rect 255 -126 317 -114
<< pdiffc >>
rect -305 -114 -271 114
rect -209 -114 -175 114
rect -113 -114 -79 114
rect -17 -114 17 114
rect 79 -114 113 114
rect 175 -114 209 114
rect 271 -114 305 114
<< poly >>
rect -177 207 -111 223
rect -177 173 -161 207
rect -127 173 -111 207
rect -177 157 -111 173
rect 15 207 81 223
rect 15 173 31 207
rect 65 173 81 207
rect 15 157 81 173
rect 207 207 273 223
rect 207 173 223 207
rect 257 173 273 207
rect 207 157 273 173
rect -255 126 -225 152
rect -159 126 -129 157
rect -63 126 -33 152
rect 33 126 63 157
rect 129 126 159 152
rect 225 126 255 157
rect -255 -157 -225 -126
rect -159 -152 -129 -126
rect -63 -157 -33 -126
rect 33 -152 63 -126
rect 129 -157 159 -126
rect 225 -152 255 -126
rect -273 -173 -207 -157
rect -273 -207 -257 -173
rect -223 -207 -207 -173
rect -273 -223 -207 -207
rect -81 -173 -15 -157
rect -81 -207 -65 -173
rect -31 -207 -15 -173
rect -81 -223 -15 -207
rect 111 -173 177 -157
rect 111 -207 127 -173
rect 161 -207 177 -173
rect 111 -223 177 -207
<< polycont >>
rect -161 173 -127 207
rect 31 173 65 207
rect 223 173 257 207
rect -257 -207 -223 -173
rect -65 -207 -31 -173
rect 127 -207 161 -173
<< locali >>
rect -177 173 -161 207
rect -127 173 -111 207
rect 15 173 31 207
rect 65 173 81 207
rect 207 173 223 207
rect 257 173 273 207
rect -305 114 -271 130
rect -305 -130 -271 -114
rect -209 114 -175 130
rect -209 -130 -175 -114
rect -113 114 -79 130
rect -113 -130 -79 -114
rect -17 114 17 130
rect -17 -130 17 -114
rect 79 114 113 130
rect 79 -130 113 -114
rect 175 114 209 130
rect 175 -130 209 -114
rect 271 114 305 130
rect 271 -130 305 -114
rect -273 -207 -257 -173
rect -223 -207 -207 -173
rect -81 -207 -65 -173
rect -31 -207 -15 -173
rect 111 -207 127 -173
rect 161 -207 177 -173
<< viali >>
rect -305 -114 -271 114
rect -209 -114 -175 114
rect -113 -114 -79 114
rect -17 -114 17 114
rect 79 -114 113 114
rect 175 -114 209 114
rect 271 -114 305 114
<< metal1 >>
rect -311 114 -265 126
rect -311 -114 -305 114
rect -271 -114 -265 114
rect -311 -126 -265 -114
rect -215 114 -169 126
rect -215 -114 -209 114
rect -175 -114 -169 114
rect -215 -126 -169 -114
rect -119 114 -73 126
rect -119 -114 -113 114
rect -79 -114 -73 114
rect -119 -126 -73 -114
rect -23 114 23 126
rect -23 -114 -17 114
rect 17 -114 23 114
rect -23 -126 23 -114
rect 73 114 119 126
rect 73 -114 79 114
rect 113 -114 119 114
rect 73 -126 119 -114
rect 169 114 215 126
rect 169 -114 175 114
rect 209 -114 215 114
rect 169 -126 215 -114
rect 265 114 311 126
rect 265 -114 271 114
rect 305 -114 311 114
rect 265 -126 311 -114
<< properties >>
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 1.26 l 0.15 m 1 nf 6 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 0 botc 0 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 0 viasrc 100 viadrn 100 viagate 0 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
